* Multi-domian SPICE model
V1 in 0 SINE(0 2.1 1k 0 0 0 10)
Rsh 0 N0 0.00000001
B1 Q 0 V=idt(-I(Rsh))

*Grain_0:
XU_0 in N0 fe_tanh Vc=0.9777151714554085 Qo=0.11823853722601885 K=2.62 tau=0.11823853722601885

*Grain_1:
XU_1 in N0 fe_tanh Vc=1.170751650546949 Qo=0.09598743247917832 K=2.62 tau=0.09598743247917832

*Grain_2:
XU_2 in N0 fe_tanh Vc=1.0201581200960494 Qo=0.09720271745313387 K=2.62 tau=0.09720271745313387

*Grain_3:
XU_3 in N0 fe_tanh Vc=0.9577680865499073 Qo=0.09167598535718255 K=2.62 tau=0.09167598535718255

*Grain_4:
XU_4 in N0 fe_tanh Vc=0.9266496933023997 Qo=0.10527566699499193 K=2.62 tau=0.10527566699499193

*Grain_5:
XU_5 in N0 fe_tanh Vc=0.8700850309035738 Qo=0.11040658070427133 K=2.62 tau=0.11040658070427133

*Grain_6:
XU_6 in N0 fe_tanh Vc=0.8485157777719095 Qo=0.09189095019986017 K=2.62 tau=0.09189095019986017

*Grain_7:
XU_7 in N0 fe_tanh Vc=0.9759124514293696 Qo=0.10265082199990497 K=2.62 tau=0.10265082199990497

*Grain_8:
XU_8 in N0 fe_tanh Vc=1.0474195546850482 Qo=0.09282611363061506 K=2.62 tau=0.09282611363061506

*Grain_9:
XU_9 in N0 fe_tanh Vc=1.19775584160247 Qo=0.09384519395484284 K=2.62 tau=0.09384519395484284
.tran 0 1.5m 0 1e-9

.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.backanno
.end
