* Multi-domian SPICE model
V1 in 0 SINE(0 2.1 1k 0 0 0 10)
Rsh 0 N0 0.00000001
B1 Q 0 V=idt(-I(Rsh))

*Grain_0:
XU_0 in N0 fe_tanh Vc=0.8802563060278936 Qo=0.10275559046295768 K=2.62 tau=0.10275559046295768

*Grain_1:
XU_1 in N0 fe_tanh Vc=1.03302630484089 Qo=0.09851785471281012 K=2.62 tau=0.09851785471281012

*Grain_2:
XU_2 in N0 fe_tanh Vc=0.9540818203316281 Qo=0.10058921674380758 K=2.62 tau=0.10058921674380758

*Grain_3:
XU_3 in N0 fe_tanh Vc=1.0362591795002183 Qo=0.10594305307600943 K=2.62 tau=0.10594305307600943

*Grain_4:
XU_4 in N0 fe_tanh Vc=0.9634887816889046 Qo=0.08749320006197514 K=2.62 tau=0.08749320006197514

*Grain_5:
XU_5 in N0 fe_tanh Vc=1.077283467281198 Qo=0.09621645253328534 K=2.62 tau=0.09621645253328534

*Grain_6:
XU_6 in N0 fe_tanh Vc=0.8962574202319418 Qo=0.0994988147041637 K=2.62 tau=0.0994988147041637

*Grain_7:
XU_7 in N0 fe_tanh Vc=0.9563217170431716 Qo=0.09977256424423366 K=2.62 tau=0.09977256424423366

*Grain_8:
XU_8 in N0 fe_tanh Vc=1.0044411873328314 Qo=0.10900473724726953 K=2.62 tau=0.10900473724726953

*Grain_9:
XU_9 in N0 fe_tanh Vc=1.2261938303698692 Qo=0.1002085162134878 K=2.62 tau=0.1002085162134878
.tran 0 1.5m 0 1e-9

.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.backanno
.end
