* Multi-domian SPICE model
.subckt fe_tanh_md in out

*Grain_0:
XU_0 in out fe_tanh Vc=0.5106471534729239 Qo=3.805490134297339e-13 K=2.62 tau=1.0962162905768435e-07 off=-0.1

*Grain_1:
XU_1 in out fe_tanh Vc=0.034509040764962695 Qo=1.1459513068878223e-14 K=2.62 tau=9.91011316205373e-08 off=-0.1

*Grain_2:
XU_2 in out fe_tanh Vc=0.04557128991269804 Qo=1.6449478293127555e-14 K=2.62 tau=8.923007758275212e-08 off=-0.1

*Grain_3:
XU_3 in out fe_tanh Vc=0.3545316972249254 Qo=2.3681270637747964e-13 K=2.62 tau=1.0462161864070541e-07 off=-0.1

*Grain_4:
XU_4 in out fe_tanh Vc=0.6910221531192295 Qo=5.638881550703724e-13 K=2.62 tau=1.141482876358601e-07 off=-0.1

*Grain_5:
XU_5 in out fe_tanh Vc=0.7225984286917916 Qo=5.976122994880839e-13 K=2.62 tau=1.0290359761894417e-07 off=-0.1

*Grain_6:
XU_6 in out fe_tanh Vc=0.5959868335363174 Qo=4.652228907559991e-13 K=2.62 tau=1.036819869496836e-07 off=-0.1

*Grain_7:
XU_7 in out fe_tanh Vc=0.7201624086363843 Qo=5.949945572307296e-13 K=2.62 tau=9.176678706007163e-08 off=-0.1

*Grain_8:
XU_8 in out fe_tanh Vc=0.254684910184114 Qo=1.5404854081511765e-13 K=2.62 tau=1.0424457950095651e-07 off=-0.1

*Grain_9:
XU_9 in out fe_tanh Vc=0.6970744996229458 Qo=5.703170624808026e-13 K=2.62 tau=9.856287555852747e-08 off=-0.1

*Grain_10:
XU_10 in out fe_tanh Vc=0.4470904268087553 Qo=3.2016023673948897e-13 K=2.62 tau=9.964304020146299e-08 off=-0.1

*Grain_11:
XU_11 in out fe_tanh Vc=0.6720770481134002 Qo=5.438738699029444e-13 K=2.62 tau=1.0898103961690038e-07 off=-0.1

*Grain_12:
XU_12 in out fe_tanh Vc=0.6636840802412625 Qo=5.350609187113209e-13 K=2.62 tau=1.0304556030489124e-07 off=-0.1

*Grain_13:
XU_13 in out fe_tanh Vc=0.45819089588329875 Qo=3.3053222168780654e-13 K=2.62 tau=9.231104716707023e-08 off=-0.1

*Grain_14:
XU_14 in out fe_tanh Vc=0.471004108946963 Qo=3.4259854565084473e-13 K=2.62 tau=1.0857346216752861e-07 off=-0.1

*Grain_15:
XU_15 in out fe_tanh Vc=0.3381257663822988 Qo=2.2266664078716991e-13 K=2.62 tau=1.0766515518816212e-07 off=-0.1

*Grain_16:
XU_16 in out fe_tanh Vc=0.0071711871063316335 Qo=1.4863523723308907e-15 K=2.62 tau=1.2041390848709714e-07 off=-0.1

*Grain_17:
XU_17 in out fe_tanh Vc=0.6360474315490521 Qo=5.062788262992564e-13 K=2.62 tau=9.216257641479182e-08 off=-0.1

*Grain_18:
XU_18 in out fe_tanh Vc=0.2780152324171137 Qo=1.7264045796190667e-13 K=2.62 tau=9.687514163380913e-08 off=-0.1

*Grain_19:
XU_19 in out fe_tanh Vc=0.41215681862516657 Qo=2.880279585403567e-13 K=2.62 tau=1.0408635749823978e-07 off=-0.1

*Grain_20:
XU_20 in out fe_tanh Vc=0.23930535109391013 Qo=1.420664549274601e-13 K=2.62 tau=1.0554550933902753e-07 off=-0.1

*Grain_21:
XU_21 in out fe_tanh Vc=-0.30129383207809757 Qo=1.9166407781663745e-13 K=2.62 tau=9.461463435418202e-08 off=-0.1

*Grain_22:
XU_22 in out fe_tanh Vc=0.4937446574384348 Qo=3.642558561192344e-13 K=2.62 tau=1.0107537550161913e-07 off=-0.1

*Grain_23:
XU_23 in out fe_tanh Vc=0.43916762941554255 Qo=3.128043817678901e-13 K=2.62 tau=1.0068164513465239e-07 off=-0.1

*Grain_24:
XU_24 in out fe_tanh Vc=0.36738083049759446 Qo=2.4803036335041665e-13 K=2.62 tau=1.008253446087289e-07 off=-0.1

*Grain_25:
XU_25 in out fe_tanh Vc=0.38274222831361043 Qo=2.615963654482451e-13 K=2.62 tau=9.9705635140268e-08 off=-0.1

*Grain_26:
XU_26 in out fe_tanh Vc=0.5490116403697967 Qo=4.181281711288716e-13 K=2.62 tau=9.317570821684333e-08 off=-0.1

*Grain_27:
XU_27 in out fe_tanh Vc=0.05186576483463701 Qo=1.9462491368663226e-14 K=2.62 tau=1.1257801098867917e-07 off=-0.1

*Grain_28:
XU_28 in out fe_tanh Vc=0.408211939096291 Qo=2.844492700927109e-13 K=2.62 tau=1.0514642949720805e-07 off=-0.1

*Grain_29:
XU_29 in out fe_tanh Vc=0.421386109440304 Qo=2.964406047003905e-13 K=2.62 tau=9.64001545178759e-08 off=-0.1

*Grain_30:
XU_30 in out fe_tanh Vc=0.12095209105127447 Qo=5.851278987812875e-14 K=2.62 tau=1.0012621988355065e-07 off=-0.1

*Grain_31:
XU_31 in out fe_tanh Vc=0.3393409321019454 Qo=2.2370749429479878e-13 K=2.62 tau=8.816105140192096e-08 off=-0.1

*Grain_32:
XU_32 in out fe_tanh Vc=0.7478763994936585 Qo=6.249311711634962e-13 K=2.62 tau=1.116181320690554e-07 off=-0.1

*Grain_33:
XU_33 in out fe_tanh Vc=0.6657522048892317 Qo=5.37229445024262e-13 K=2.62 tau=9.257895529114622e-08 off=-0.1

*Grain_34:
XU_34 in out fe_tanh Vc=0.9017248813139058 Qo=7.969841413889351e-13 K=2.62 tau=9.14837823010427e-08 off=-0.1

*Grain_35:
XU_35 in out fe_tanh Vc=0.4720883472786169 Qo=3.436241474695101e-13 K=2.62 tau=9.195110658638605e-08 off=-0.1

*Grain_36:
XU_36 in out fe_tanh Vc=0.666421816196064 Qo=5.379319975940025e-13 K=2.62 tau=9.804889197467341e-08 off=-0.1

*Grain_37:
XU_37 in out fe_tanh Vc=0.05003088982747039 Qo=1.8572189473609665e-14 K=2.62 tau=1.0640903148106343e-07 off=-0.1

*Grain_38:
XU_38 in out fe_tanh Vc=0.8923700711311644 Qo=7.862522576852245e-13 K=2.62 tau=1.016281533436246e-07 off=-0.1

*Grain_39:
XU_39 in out fe_tanh Vc=0.8737171443397338 Qo=7.649543618743388e-13 K=2.62 tau=1.0743320796084023e-07 off=-0.1

*Grain_40:
XU_40 in out fe_tanh Vc=0.43740460423298233 Qo=3.1117289884917385e-13 K=2.62 tau=1.031638649828301e-07 off=-0.1

*Grain_41:
XU_41 in out fe_tanh Vc=-0.15494297277402924 Qo=8.073779044534385e-14 K=2.62 tau=8.842422459432844e-08 off=-0.1

*Grain_42:
XU_42 in out fe_tanh Vc=0.21218677617224016 Qo=1.2150306102177873e-13 K=2.62 tau=1.100408544332784e-07 off=-0.1

*Grain_43:
XU_43 in out fe_tanh Vc=-0.03244478511327947 Qo=1.0576495359169422e-14 K=2.62 tau=7.399959160493193e-08 off=-0.1

*Grain_44:
XU_44 in out fe_tanh Vc=0.017347890324461934 Qo=4.686774718753001e-15 K=2.62 tau=9.791343613337152e-08 off=-0.1

*Grain_45:
XU_45 in out fe_tanh Vc=0.2724547395409157 Qo=1.6816518435972167e-13 K=2.62 tau=1.0145021739416984e-07 off=-0.1

*Grain_46:
XU_46 in out fe_tanh Vc=0.7019020654285337 Qo=5.75457012753123e-13 K=2.62 tau=9.594325678713977e-08 off=-0.1

*Grain_47:
XU_47 in out fe_tanh Vc=0.5124398670614696 Qo=3.822867038234443e-13 K=2.62 tau=9.396458462281162e-08 off=-0.1

*Grain_48:
XU_48 in out fe_tanh Vc=-0.450991490552784 Qo=3.2379658365911854e-13 K=2.62 tau=1.1669820137539725e-07 off=-0.1

*Grain_49:
XU_49 in out fe_tanh Vc=0.22556869902261673 Qo=1.315575859224852e-13 K=2.62 tau=9.871523411867602e-08 off=-0.1

*Grain_50:
XU_50 in out fe_tanh Vc=0.1819111425916337 Qo=9.946504939229334e-14 K=2.62 tau=8.30460839358074e-08 off=-0.1

*Grain_51:
XU_51 in out fe_tanh Vc=0.7704018513606201 Qo=6.495101220145994e-13 K=2.62 tau=9.048598686956934e-08 off=-0.1

*Grain_52:
XU_52 in out fe_tanh Vc=0.3805813910427512 Qo=2.596780398830814e-13 K=2.62 tau=1.0674961482899544e-07 off=-0.1

*Grain_53:
XU_53 in out fe_tanh Vc=0.7142840527825952 Qo=5.886886339180354e-13 K=2.62 tau=1.0588734945573379e-07 off=-0.1

*Grain_54:
XU_54 in out fe_tanh Vc=0.4566419164438684 Qo=3.2908032440151295e-13 K=2.62 tau=1.0629318962561583e-07 off=-0.1

*Grain_55:
XU_55 in out fe_tanh Vc=0.3310621965040311 Qo=2.1663861984505103e-13 K=2.62 tau=1.0753997045451263e-07 off=-0.1

*Grain_56:
XU_56 in out fe_tanh Vc=0.3818755147649882 Qo=2.608265322394648e-13 K=2.62 tau=1.108091839825998e-07 off=-0.1

*Grain_57:
XU_57 in out fe_tanh Vc=0.5784557981917602 Qo=4.47511955945116e-13 K=2.62 tau=9.912137858866086e-08 off=-0.1

*Grain_58:
XU_58 in out fe_tanh Vc=-0.025089136780016175 Qo=7.571550884549433e-15 K=2.62 tau=8.895690858320637e-08 off=-0.1

*Grain_59:
XU_59 in out fe_tanh Vc=0.5098087742035972 Qo=3.7973699373911815e-13 K=2.62 tau=9.661849955937383e-08 off=-0.1

*Grain_60:
XU_60 in out fe_tanh Vc=0.1424608419136431 Qo=7.23864984494252e-14 K=2.62 tau=1.1706082869245841e-07 off=-0.1

*Grain_61:
XU_61 in out fe_tanh Vc=0.0612718974280535 Qo=2.417091765196076e-14 K=2.62 tau=1.0824697547045302e-07 off=-0.1

*Grain_62:
XU_62 in out fe_tanh Vc=0.21740328355840766 Qo=1.2540052057047733e-13 K=2.62 tau=1.0680771903477749e-07 off=-0.1

*Grain_63:
XU_63 in out fe_tanh Vc=0.2378587353431391 Qo=1.409510279642261e-13 K=2.62 tau=1.0146103672492908e-07 off=-0.1

*Grain_64:
XU_64 in out fe_tanh Vc=0.321699201795904 Qo=2.0870765995108585e-13 K=2.62 tau=8.658225473720289e-08 off=-0.1

*Grain_65:
XU_65 in out fe_tanh Vc=0.6431515834082223 Qo=5.136422699298911e-13 K=2.62 tau=1.0265531072371162e-07 off=-0.1

*Grain_66:
XU_66 in out fe_tanh Vc=0.00247966737237576 Qo=3.7373594247647703e-16 K=2.62 tau=1.1320510271091626e-07 off=-0.1

*Grain_67:
XU_67 in out fe_tanh Vc=0.8225184717156263 Qo=7.072008407396604e-13 K=2.62 tau=1.1203364106599983e-07 off=-0.1

*Grain_68:
XU_68 in out fe_tanh Vc=0.5765250764220655 Qo=4.4557116010410524e-13 K=2.62 tau=9.376664129811582e-08 off=-0.1

*Grain_69:
XU_69 in out fe_tanh Vc=-0.1481856371461897 Qo=7.619059335597101e-14 K=2.62 tau=1.0455685901786864e-07 off=-0.1

*Grain_70:
XU_70 in out fe_tanh Vc=0.17727512716107424 Qo=9.618238848980472e-14 K=2.62 tau=1.0540440911680003e-07 off=-0.1

*Grain_71:
XU_71 in out fe_tanh Vc=0.5067060961067853 Qo=3.7673535471405506e-13 K=2.62 tau=1.0116164659801462e-07 off=-0.1

*Grain_72:
XU_72 in out fe_tanh Vc=0.7938945597127962 Qo=6.753751610050384e-13 K=2.62 tau=1.0047345052059981e-07 off=-0.1

*Grain_73:
XU_73 in out fe_tanh Vc=0.47675346461988927 Qo=3.480450212215951e-13 K=2.62 tau=1.0139377560259903e-07 off=-0.1

*Grain_74:
XU_74 in out fe_tanh Vc=0.4736722729126591 Qo=3.4512368340169357e-13 K=2.62 tau=1.0245099081328611e-07 off=-0.1

*Grain_75:
XU_75 in out fe_tanh Vc=0.5415703600366594 Qo=4.107757187564698e-13 K=2.62 tau=9.65312200888537e-08 off=-0.1

*Grain_76:
XU_76 in out fe_tanh Vc=0.942425841819516 Qo=8.440627849497723e-13 K=2.62 tau=8.172452797172458e-08 off=-0.1

*Grain_77:
XU_77 in out fe_tanh Vc=0.43503756840059254 Qo=3.089855730284756e-13 K=2.62 tau=9.74552729855123e-08 off=-0.1

*Grain_78:
XU_78 in out fe_tanh Vc=-0.04527334979351394 Qo=1.630980724900958e-14 K=2.62 tau=9.251894974794175e-08 off=-0.1

*Grain_79:
XU_79 in out fe_tanh Vc=0.13070275680421162 Qo=6.47177757286249e-14 K=2.62 tau=1.0571172131179094e-07 off=-0.1

*Grain_80:
XU_80 in out fe_tanh Vc=0.28534112617609386 Qo=1.7857764553593314e-13 K=2.62 tau=9.869243615384484e-08 off=-0.1

*Grain_81:
XU_81 in out fe_tanh Vc=-0.19079366045591006 Qo=1.0582457493000495e-13 K=2.62 tau=1.0509717842041741e-07 off=-0.1

*Grain_82:
XU_82 in out fe_tanh Vc=0.2558906173522638 Qo=1.5499728149067098e-13 K=2.62 tau=1.0588946278455361e-07 off=-0.1

*Grain_83:
XU_83 in out fe_tanh Vc=-0.010946958316894961 Qo=2.5759350838234927e-15 K=2.62 tau=1.0794306720460618e-07 off=-0.1

*Grain_84:
XU_84 in out fe_tanh Vc=0.6347721648626482 Qo=5.049596162999336e-13 K=2.62 tau=9.446563270059917e-08 off=-0.1

*Grain_85:
XU_85 in out fe_tanh Vc=0.5656499510859071 Qo=4.3467582844138264e-13 K=2.62 tau=1.0768163137066455e-07 off=-0.1

*Grain_86:
XU_86 in out fe_tanh Vc=0.13622668202326127 Qo=6.829583875616517e-14 K=2.62 tau=1.0288828652555213e-07 off=-0.1

*Grain_87:
XU_87 in out fe_tanh Vc=0.9350634662375953 Qo=8.355007156092995e-13 K=2.62 tau=1.1357601102961895e-07 off=-0.1

*Grain_88:
XU_88 in out fe_tanh Vc=0.6916807357649317 Qo=5.645868968378467e-13 K=2.62 tau=1.1183391442234295e-07 off=-0.1

*Grain_89:
XU_89 in out fe_tanh Vc=0.4983282157551743 Qo=3.686578889093163e-13 K=2.62 tau=9.295220630550605e-08 off=-0.1

*Grain_90:
XU_90 in out fe_tanh Vc=0.4914898768853065 Qo=3.6209486066760153e-13 K=2.62 tau=1.1815182736774631e-07 off=-0.1

*Grain_91:
XU_91 in out fe_tanh Vc=-0.025487593339758696 Qo=7.728245122246246e-15 K=2.62 tau=1.0140795083875405e-07 off=-0.1

*Grain_92:
XU_92 in out fe_tanh Vc=0.447221906168929 Qo=3.2028263975344404e-13 K=2.62 tau=1.21432463129927e-07 off=-0.1

*Grain_93:
XU_93 in out fe_tanh Vc=0.3945797302305776 Qo=2.7216270546791403e-13 K=2.62 tau=9.030667424451035e-08 off=-0.1

*Grain_94:
XU_94 in out fe_tanh Vc=-0.19030779768582096 Qo=1.0547437702442191e-13 K=2.62 tau=8.265864604792056e-08 off=-0.1

*Grain_95:
XU_95 in out fe_tanh Vc=0.6852459108473695 Qo=5.577682623885562e-13 K=2.62 tau=1.072321340592539e-07 off=-0.1

*Grain_96:
XU_96 in out fe_tanh Vc=0.4523552673089687 Qo=3.250700496776519e-13 K=2.62 tau=9.015241398475668e-08 off=-0.1

*Grain_97:
XU_97 in out fe_tanh Vc=0.5857621838135446 Qo=4.548740277037931e-13 K=2.62 tau=1.0908597866655548e-07 off=-0.1

*Grain_98:
XU_98 in out fe_tanh Vc=0.896910909294607 Qo=7.914573358249748e-13 K=2.62 tau=8.943076645010305e-08 off=-0.1

*Grain_99:
XU_99 in out fe_tanh Vc=0.5597103703427955 Qo=4.287516161796279e-13 K=2.62 tau=1.0655768638275021e-07 off=-0.1

*Grain_100:
XU_100 in out fe_tanh Vc=0.33899805592511967 Qo=2.2341368934706832e-13 K=2.62 tau=1.1139282399816895e-07 off=-0.1

*Grain_101:
XU_101 in out fe_tanh Vc=0.7000423107591036 Qo=5.734756562259294e-13 K=2.62 tau=1.0723246595777235e-07 off=-0.1

*Grain_102:
XU_102 in out fe_tanh Vc=0.8102748788655899 Qo=6.935463610641415e-13 K=2.62 tau=1.0213578673307348e-07 off=-0.1

*Grain_103:
XU_103 in out fe_tanh Vc=0.5930916056195481 Qo=4.62287042646334e-13 K=2.62 tau=1.0368185718280751e-07 off=-0.1

*Grain_104:
XU_104 in out fe_tanh Vc=0.8951268840463815 Qo=7.894113958182006e-13 K=2.62 tau=1.0136879801484785e-07 off=-0.1

*Grain_105:
XU_105 in out fe_tanh Vc=0.4679276426726038 Qo=3.3969231574750903e-13 K=2.62 tau=1.0928865928363543e-07 off=-0.1

*Grain_106:
XU_106 in out fe_tanh Vc=0.43474363877765904 Qo=3.087142078453302e-13 K=2.62 tau=9.384740543063667e-08 off=-0.1

*Grain_107:
XU_107 in out fe_tanh Vc=0.24884510414934696 Qo=1.4947248038620055e-13 K=2.62 tau=1.0258270195035354e-07 off=-0.1

*Grain_108:
XU_108 in out fe_tanh Vc=0.18006433362389854 Qo=9.815431985146824e-14 K=2.62 tau=1.0091435131168373e-07 off=-0.1

*Grain_109:
XU_109 in out fe_tanh Vc=0.4206961733938076 Qo=2.9580978833964235e-13 K=2.62 tau=1.0689565381549604e-07 off=-0.1

*Grain_110:
XU_110 in out fe_tanh Vc=0.7291586732901989 Qo=6.046750794104524e-13 K=2.62 tau=9.756889073612524e-08 off=-0.1

*Grain_111:
XU_111 in out fe_tanh Vc=-0.0902028794157701 Qo=3.99613297997327e-14 K=2.62 tau=1.2048320267199017e-07 off=-0.1

*Grain_112:
XU_112 in out fe_tanh Vc=0.3628930630824013 Qo=2.4409881823619206e-13 K=2.62 tau=1.1063044937997449e-07 off=-0.1

*Grain_113:
XU_113 in out fe_tanh Vc=-0.10249229103330793 Qo=4.717935202801642e-14 K=2.62 tau=1.170366741381858e-07 off=-0.1

*Grain_114:
XU_114 in out fe_tanh Vc=0.6078628223901854 Qo=4.77310147359191e-13 K=2.62 tau=1.0000206661769974e-07 off=-0.1

*Grain_115:
XU_115 in out fe_tanh Vc=0.5017609673922581 Qo=3.719626615524179e-13 K=2.62 tau=9.720301719966569e-08 off=-0.1

*Grain_116:
XU_116 in out fe_tanh Vc=0.5308386431715857 Qo=4.0022544853203876e-13 K=2.62 tau=6.63149769393353e-08 off=-0.1

*Grain_117:
XU_117 in out fe_tanh Vc=0.17589162566890157 Qo=9.520771061802193e-14 K=2.62 tau=1.1441278831850239e-07 off=-0.1

*Grain_118:
XU_118 in out fe_tanh Vc=0.757938432108358 Qo=6.358834445802485e-13 K=2.62 tau=9.720126777193424e-08 off=-0.1

*Grain_119:
XU_119 in out fe_tanh Vc=0.41921620738313886 Qo=2.9445768572337126e-13 K=2.62 tau=1.00828856452347e-07 off=-0.1

*Grain_120:
XU_120 in out fe_tanh Vc=0.5047180714031426 Qo=3.748149645184187e-13 K=2.62 tau=9.5536305082145e-08 off=-0.1

*Grain_121:
XU_121 in out fe_tanh Vc=0.5401974711571186 Qo=4.09422514529971e-13 K=2.62 tau=8.587136554389206e-08 off=-0.1

*Grain_122:
XU_122 in out fe_tanh Vc=0.009397216326906543 Qo=2.1122844522594488e-15 K=2.62 tau=1.0127253167949334e-07 off=-0.1

*Grain_123:
XU_123 in out fe_tanh Vc=-0.010358219895379217 Qo=2.3973093256382256e-15 K=2.62 tau=9.112243697979203e-08 off=-0.1

*Grain_124:
XU_124 in out fe_tanh Vc=0.4885899403945707 Qo=3.593199145695662e-13 K=2.62 tau=8.711890381079436e-08 off=-0.1

*Grain_125:
XU_125 in out fe_tanh Vc=1.021907254157846 Qo=9.377527299304386e-13 K=2.62 tau=9.949579327041094e-08 off=-0.1

*Grain_126:
XU_126 in out fe_tanh Vc=0.7216237533049167 Qo=5.965645970378946e-13 K=2.62 tau=1.1303395686668656e-07 off=-0.1

*Grain_127:
XU_127 in out fe_tanh Vc=0.4205573239823073 Qo=2.9568287424038233e-13 K=2.62 tau=1.1010076822553705e-07 off=-0.1

*Grain_128:
XU_128 in out fe_tanh Vc=0.6884135163473615 Qo=5.611224124828828e-13 K=2.62 tau=1.054251670218883e-07 off=-0.1

*Grain_129:
XU_129 in out fe_tanh Vc=0.1815899094824964 Qo=9.923677365456706e-14 K=2.62 tau=9.790821738166778e-08 off=-0.1

*Grain_130:
XU_130 in out fe_tanh Vc=0.5073124758960514 Qo=3.7732155530127204e-13 K=2.62 tau=1.0158800512554376e-07 off=-0.1

*Grain_131:
XU_131 in out fe_tanh Vc=0.17888922832694848 Qo=9.732241077006769e-14 K=2.62 tau=9.630744980021036e-08 off=-0.1

*Grain_132:
XU_132 in out fe_tanh Vc=0.08920538104884596 Qo=3.938780497865969e-14 K=2.62 tau=1.1768102870666249e-07 off=-0.1

*Grain_133:
XU_133 in out fe_tanh Vc=0.8363264765178651 Qo=7.226733010960937e-13 K=2.62 tau=8.776114504558955e-08 off=-0.1

*Grain_134:
XU_134 in out fe_tanh Vc=0.13699398133749663 Qo=6.879634156217595e-14 K=2.62 tau=1.0523092700221374e-07 off=-0.1

*Grain_135:
XU_135 in out fe_tanh Vc=-0.09297057779739942 Qo=4.1562589656314466e-14 K=2.62 tau=1.0288810230554641e-07 off=-0.1

*Grain_136:
XU_136 in out fe_tanh Vc=0.42972165214000174 Qo=3.0408627474786606e-13 K=2.62 tau=9.152237508581679e-08 off=-0.1

*Grain_137:
XU_137 in out fe_tanh Vc=0.3863088353654607 Qo=2.6476979786804105e-13 K=2.62 tau=8.811710350765278e-08 off=-0.1

*Grain_138:
XU_138 in out fe_tanh Vc=0.059296634476322385 Qo=2.3162875265165097e-14 K=2.62 tau=1.0895194145460112e-07 off=-0.1

*Grain_139:
XU_139 in out fe_tanh Vc=-0.024035841434501937 Qo=7.160948325628817e-15 K=2.62 tau=8.719963362499665e-08 off=-0.1

*Grain_140:
XU_140 in out fe_tanh Vc=0.5083230787710873 Qo=3.782989942646335e-13 K=2.62 tau=9.751611789479793e-08 off=-0.1

*Grain_141:
XU_141 in out fe_tanh Vc=0.31767774606612387 Qo=2.0532235694331725e-13 K=2.62 tau=9.767264114623967e-08 off=-0.1

*Grain_142:
XU_142 in out fe_tanh Vc=0.401912589165152 Qo=2.787561792510223e-13 K=2.62 tau=9.814837585478562e-08 off=-0.1

*Grain_143:
XU_143 in out fe_tanh Vc=0.5674182575954564 Qo=4.364431765074826e-13 K=2.62 tau=1.0621745606459102e-07 off=-0.1

*Grain_144:
XU_144 in out fe_tanh Vc=0.7840501086859011 Qo=6.64508247599518e-13 K=2.62 tau=1.0186100905519949e-07 off=-0.1

*Grain_145:
XU_145 in out fe_tanh Vc=0.9758340816264032 Qo=8.831656864254698e-13 K=2.62 tau=9.131868177869574e-08 off=-0.1

*Grain_146:
XU_146 in out fe_tanh Vc=0.19173629568578707 Qo=1.0650476607515348e-13 K=2.62 tau=9.884844939052234e-08 off=-0.1

*Grain_147:
XU_147 in out fe_tanh Vc=-0.17677362352724624 Qo=9.582881415122571e-14 K=2.62 tau=1.0710087660920742e-07 off=-0.1

*Grain_148:
XU_148 in out fe_tanh Vc=0.07430816791835787 Qo=3.105996273998303e-14 K=2.62 tau=9.951451101812727e-08 off=-0.1

*Grain_149:
XU_149 in out fe_tanh Vc=0.47029477300927974 Qo=3.4192795424748487e-13 K=2.62 tau=1.0464775831117123e-07 off=-0.1

*Grain_150:
XU_150 in out fe_tanh Vc=0.4200148723171625 Qo=2.9518717151052133e-13 K=2.62 tau=1.044707171887752e-07 off=-0.1

*Grain_151:
XU_151 in out fe_tanh Vc=0.6085128566346925 Qo=4.779738053294332e-13 K=2.62 tau=9.424725665861305e-08 off=-0.1

*Grain_152:
XU_152 in out fe_tanh Vc=0.5544358620847788 Qo=4.2350653687790247e-13 K=2.62 tau=1.1527229293393959e-07 off=-0.1

*Grain_153:
XU_153 in out fe_tanh Vc=0.09370602834396019 Qo=4.1990514964541e-14 K=2.62 tau=9.143366949046981e-08 off=-0.1

*Grain_154:
XU_154 in out fe_tanh Vc=0.26484357859112906 Qo=1.6208383065115738e-13 K=2.62 tau=9.81943419531141e-08 off=-0.1

*Grain_155:
XU_155 in out fe_tanh Vc=0.30983308128557374 Qo=1.987556725241189e-13 K=2.62 tau=1.0016318162276431e-07 off=-0.1

*Grain_156:
XU_156 in out fe_tanh Vc=0.5019915719778308 Qo=3.7218491253993615e-13 K=2.62 tau=1.062285755326906e-07 off=-0.1

*Grain_157:
XU_157 in out fe_tanh Vc=0.27278656178358407 Qo=1.6843148356866535e-13 K=2.62 tau=1.1439792508644937e-07 off=-0.1

*Grain_158:
XU_158 in out fe_tanh Vc=0.855513030637882 Qo=7.443000152823722e-13 K=2.62 tau=1.0043562383178701e-07 off=-0.1

*Grain_159:
XU_159 in out fe_tanh Vc=0.656544367455827 Qo=5.275901930798566e-13 K=2.62 tau=9.149648603807583e-08 off=-0.1

*Grain_160:
XU_160 in out fe_tanh Vc=0.38970127188217046 Qo=2.677964284518423e-13 K=2.62 tau=7.974306919700541e-08 off=-0.1

*Grain_161:
XU_161 in out fe_tanh Vc=0.1371338188469765 Qo=6.888764715170475e-14 K=2.62 tau=1.1409700234648272e-07 off=-0.1

*Grain_162:
XU_162 in out fe_tanh Vc=0.359810586574477 Qo=2.414068164895271e-13 K=2.62 tau=1.0441111536967083e-07 off=-0.1

*Grain_163:
XU_163 in out fe_tanh Vc=0.3045934404986714 Qo=1.9439725172001643e-13 K=2.62 tau=8.061679289117395e-08 off=-0.1

*Grain_164:
XU_164 in out fe_tanh Vc=0.19959504802326444 Qo=1.1221427328966434e-13 K=2.62 tau=9.602795704832882e-08 off=-0.1

*Grain_165:
XU_165 in out fe_tanh Vc=0.7228861765344825 Qo=5.979216877843816e-13 K=2.62 tau=1.1198620472288942e-07 off=-0.1

*Grain_166:
XU_166 in out fe_tanh Vc=0.5431046213794501 Qo=4.122891997215662e-13 K=2.62 tau=1.0093160754202054e-07 off=-0.1

*Grain_167:
XU_167 in out fe_tanh Vc=-0.29327268992857014 Qo=1.850574271150648e-13 K=2.62 tau=9.474026355825484e-08 off=-0.1

*Grain_168:
XU_168 in out fe_tanh Vc=0.3818844880233112 Qo=2.6083449979332246e-13 K=2.62 tau=9.522382286510128e-08 off=-0.1

*Grain_169:
XU_169 in out fe_tanh Vc=-0.037547952948952745 Qo=1.2788380656237671e-14 K=2.62 tau=1.1077650556198445e-07 off=-0.1

*Grain_170:
XU_170 in out fe_tanh Vc=0.48473266327233944 Qo=3.5563654403575365e-13 K=2.62 tau=8.544724903421793e-08 off=-0.1

*Grain_171:
XU_171 in out fe_tanh Vc=0.023346804351490336 Qo=6.895235243267258e-15 K=2.62 tau=1.1176112228321882e-07 off=-0.1

*Grain_172:
XU_172 in out fe_tanh Vc=0.36617488256667385 Qo=2.4697245946832445e-13 K=2.62 tau=1.0261852949811092e-07 off=-0.1

*Grain_173:
XU_173 in out fe_tanh Vc=0.9422872097298816 Qo=8.439013769316881e-13 K=2.62 tau=1.0541525766772923e-07 off=-0.1

*Grain_174:
XU_174 in out fe_tanh Vc=-0.27977781678520686 Qo=1.740646857526942e-13 K=2.62 tau=1.194847147348393e-07 off=-0.1

*Grain_175:
XU_175 in out fe_tanh Vc=0.5088363494722202 Qo=3.787956448402421e-13 K=2.62 tau=1.1189014310305518e-07 off=-0.1

*Grain_176:
XU_176 in out fe_tanh Vc=0.46228607053071374 Qo=3.343778186733792e-13 K=2.62 tau=1.044821793721905e-07 off=-0.1

*Grain_177:
XU_177 in out fe_tanh Vc=0.24396703426665994 Qo=1.4567462248568032e-13 K=2.62 tau=1.0036982511382698e-07 off=-0.1

*Grain_178:
XU_178 in out fe_tanh Vc=0.5140818048558218 Qo=3.8387984719718563e-13 K=2.62 tau=8.47883020484051e-08 off=-0.1

*Grain_179:
XU_179 in out fe_tanh Vc=0.0899687003865195 Qo=3.982651374128977e-14 K=2.62 tau=9.063032802206571e-08 off=-0.1

*Grain_180:
XU_180 in out fe_tanh Vc=0.5442274006460903 Qo=4.133975850938129e-13 K=2.62 tau=9.540822361682133e-08 off=-0.1

*Grain_181:
XU_181 in out fe_tanh Vc=0.7207468034410154 Qo=5.956223048773381e-13 K=2.62 tau=8.718236969106514e-08 off=-0.1

*Grain_182:
XU_182 in out fe_tanh Vc=0.517784598995164 Qo=3.874782036124355e-13 K=2.62 tau=9.192117846439834e-08 off=-0.1

*Grain_183:
XU_183 in out fe_tanh Vc=0.253899602766394 Qo=1.5343132596467792e-13 K=2.62 tau=1.1414174043999512e-07 off=-0.1

*Grain_184:
XU_184 in out fe_tanh Vc=0.7849370992750797 Qo=6.654856931907745e-13 K=2.62 tau=9.227853755093313e-08 off=-0.1

*Grain_185:
XU_185 in out fe_tanh Vc=0.26434363701788705 Qo=1.6168619088830023e-13 K=2.62 tau=1.0607752966817709e-07 off=-0.1

*Grain_186:
XU_186 in out fe_tanh Vc=0.5327117352838001 Qo=4.020623009819454e-13 K=2.62 tau=1.0754236908074748e-07 off=-0.1

*Grain_187:
XU_187 in out fe_tanh Vc=0.6778788769919258 Qo=5.499853763676185e-13 K=2.62 tau=1.1885807414670222e-07 off=-0.1

*Grain_188:
XU_188 in out fe_tanh Vc=0.34029306425255246 Qo=2.2452382755756622e-13 K=2.62 tau=9.779988930723657e-08 off=-0.1

*Grain_189:
XU_189 in out fe_tanh Vc=0.5196508167877841 Qo=3.8929471599011855e-13 K=2.62 tau=9.228981166626394e-08 off=-0.1

*Grain_190:
XU_190 in out fe_tanh Vc=0.28144776385797166 Qo=1.754165453036394e-13 K=2.62 tau=8.709201859462091e-08 off=-0.1

*Grain_191:
XU_191 in out fe_tanh Vc=0.9736270644740651 Qo=8.805699067472741e-13 K=2.62 tau=9.804624086840182e-08 off=-0.1

*Grain_192:
XU_192 in out fe_tanh Vc=0.6558301261978827 Qo=5.268441738412314e-13 K=2.62 tau=8.650153633985384e-08 off=-0.1

*Grain_193:
XU_193 in out fe_tanh Vc=0.6487261671953779 Qo=5.194374422459438e-13 K=2.62 tau=8.473407387185205e-08 off=-0.1

*Grain_194:
XU_194 in out fe_tanh Vc=0.29201625767858885 Qo=1.8402742559358731e-13 K=2.62 tau=8.807363334611642e-08 off=-0.1

*Grain_195:
XU_195 in out fe_tanh Vc=0.25769701894808705 Qo=1.5642120366213937e-13 K=2.62 tau=1.037620887518694e-07 off=-0.1

*Grain_196:
XU_196 in out fe_tanh Vc=-0.38499231813851853 Qo=2.635973826139327e-13 K=2.62 tau=1.0805290614195228e-07 off=-0.1

*Grain_197:
XU_197 in out fe_tanh Vc=-0.026310183776539542 Qo=8.05405250658713e-15 K=2.62 tau=8.813041999646287e-08 off=-0.1

*Grain_198:
XU_198 in out fe_tanh Vc=0.28373616028542104 Qo=1.7727296307002877e-13 K=2.62 tau=9.579890064845068e-08 off=-0.1

*Grain_199:
XU_199 in out fe_tanh Vc=-0.2706855046348645 Qo=1.6674695426480347e-13 K=2.62 tau=1.0114782177246584e-07 off=-0.1

*Grain_200:
XU_200 in out fe_tanh Vc=0.4929538765781798 Qo=3.6349762911379947e-13 K=2.62 tau=1.047101561133019e-07 off=-0.1

*Grain_201:
XU_201 in out fe_tanh Vc=0.44917246044326925 Qo=3.220998093700696e-13 K=2.62 tau=9.887567109220483e-08 off=-0.1

*Grain_202:
XU_202 in out fe_tanh Vc=0.4970982045975095 Qo=3.6747539328895963e-13 K=2.62 tau=9.631564746621201e-08 off=-0.1

*Grain_203:
XU_203 in out fe_tanh Vc=0.4481903379853805 Qo=3.211845507955338e-13 K=2.62 tau=1.0977948058846203e-07 off=-0.1

*Grain_204:
XU_204 in out fe_tanh Vc=0.41289113973263913 Qo=2.886952530045671e-13 K=2.62 tau=1.1109404795466857e-07 off=-0.1

*Grain_205:
XU_205 in out fe_tanh Vc=0.3484095648813857 Qo=2.3151039734820695e-13 K=2.62 tau=1.0555430676158576e-07 off=-0.1

*Grain_206:
XU_206 in out fe_tanh Vc=0.6140805860112095 Qo=4.83666923328444e-13 K=2.62 tau=1.085948788133416e-07 off=-0.1

*Grain_207:
XU_207 in out fe_tanh Vc=0.5240654070467572 Qo=3.935995124615797e-13 K=2.62 tau=9.621111587624429e-08 off=-0.1

*Grain_208:
XU_208 in out fe_tanh Vc=0.4253560207890842 Qo=3.0007635115528837e-13 K=2.62 tau=8.461182461581119e-08 off=-0.1

*Grain_209:
XU_209 in out fe_tanh Vc=0.7852038345162287 Qo=6.657796948307551e-13 K=2.62 tau=9.54643304655641e-08 off=-0.1

*Grain_210:
XU_210 in out fe_tanh Vc=0.8486704711507211 Qo=7.365703443114863e-13 K=2.62 tau=9.069431067836036e-08 off=-0.1

*Grain_211:
XU_211 in out fe_tanh Vc=0.02583569728718249 Qo=7.865741216283863e-15 K=2.62 tau=9.553191453828093e-08 off=-0.1

*Grain_212:
XU_212 in out fe_tanh Vc=0.3386348410759195 Qo=2.231025537515646e-13 K=2.62 tau=9.514965327003724e-08 off=-0.1

*Grain_213:
XU_213 in out fe_tanh Vc=0.6168706392949931 Qo=4.865256487048921e-13 K=2.62 tau=8.571955168225982e-08 off=-0.1

*Grain_214:
XU_214 in out fe_tanh Vc=0.6281816111923779 Qo=4.981546576919883e-13 K=2.62 tau=1.033563566615005e-07 off=-0.1

*Grain_215:
XU_215 in out fe_tanh Vc=0.8354598097299548 Qo=7.216998948213066e-13 K=2.62 tau=9.932645127241843e-08 off=-0.1

*Grain_216:
XU_216 in out fe_tanh Vc=1.0633229618003655 Qo=9.874569262954932e-13 K=2.62 tau=8.107120531819779e-08 off=-0.1

*Grain_217:
XU_217 in out fe_tanh Vc=-0.15629107995784175 Qo=8.165219427064189e-14 K=2.62 tau=9.062802982488712e-08 off=-0.1

*Grain_218:
XU_218 in out fe_tanh Vc=-0.08741255886002608 Qo=3.836183687121491e-14 K=2.62 tau=1.0624826758459865e-07 off=-0.1

*Grain_219:
XU_219 in out fe_tanh Vc=0.15991177579525917 Qo=8.411975329626834e-14 K=2.62 tau=1.0662770918442137e-07 off=-0.1

*Grain_220:
XU_220 in out fe_tanh Vc=0.6134362088704334 Qo=4.830072390742379e-13 K=2.62 tau=9.698816178569104e-08 off=-0.1

*Grain_221:
XU_221 in out fe_tanh Vc=0.27617391102477223 Qo=1.7115549849594955e-13 K=2.62 tau=9.89290698467915e-08 off=-0.1

*Grain_222:
XU_222 in out fe_tanh Vc=0.04898194994697369 Qo=1.8067593116854726e-14 K=2.62 tau=1.0279298753232953e-07 off=-0.1

*Grain_223:
XU_223 in out fe_tanh Vc=0.4662696635699986 Qo=3.3812845401840127e-13 K=2.62 tau=1.0846474406672518e-07 off=-0.1

*Grain_224:
XU_224 in out fe_tanh Vc=0.44460023273890076 Qo=3.1784398848374157e-13 K=2.62 tau=9.810908545160303e-08 off=-0.1

*Grain_225:
XU_225 in out fe_tanh Vc=0.06626800962535356 Qo=2.676384555699674e-14 K=2.62 tau=8.97642422701823e-08 off=-0.1

*Grain_226:
XU_226 in out fe_tanh Vc=0.5092952061363023 Qo=3.792397706106021e-13 K=2.62 tau=1.0780827898050661e-07 off=-0.1

*Grain_227:
XU_227 in out fe_tanh Vc=0.5139288931487415 Qo=3.837314151112536e-13 K=2.62 tau=1.0805273522854272e-07 off=-0.1

*Grain_228:
XU_228 in out fe_tanh Vc=-0.22905555666631428 Qo=1.3420740893714674e-13 K=2.62 tau=1.1122784181720403e-07 off=-0.1

*Grain_229:
XU_229 in out fe_tanh Vc=0.13262951958044306 Qo=6.596076226844074e-14 K=2.62 tau=1.0912806116002782e-07 off=-0.1

*Grain_230:
XU_230 in out fe_tanh Vc=0.6816466709108517 Qo=5.539627006355026e-13 K=2.62 tau=9.370834675429117e-08 off=-0.1

*Grain_231:
XU_231 in out fe_tanh Vc=0.3810698294873726 Qo=2.601113755537577e-13 K=2.62 tau=1.0491881448404672e-07 off=-0.1

*Grain_232:
XU_232 in out fe_tanh Vc=0.12294523651762523 Qo=5.976936326505425e-14 K=2.62 tau=1.0535851126244598e-07 off=-0.1

*Grain_233:
XU_233 in out fe_tanh Vc=0.09202273735395788 Qo=4.101258114367712e-14 K=2.62 tau=9.384413499429682e-08 off=-0.1

*Grain_234:
XU_234 in out fe_tanh Vc=0.32464924988490695 Qo=2.1119913508311874e-13 K=2.62 tau=9.112428977703288e-08 off=-0.1

*Grain_235:
XU_235 in out fe_tanh Vc=0.46630311085933374 Qo=3.3815998616309835e-13 K=2.62 tau=9.556161362714659e-08 off=-0.1

*Grain_236:
XU_236 in out fe_tanh Vc=0.6035758935251156 Qo=4.729387097382379e-13 K=2.62 tau=1.0830730132728314e-07 off=-0.1

*Grain_237:
XU_237 in out fe_tanh Vc=0.2410797294484722 Qo=1.4343737028270033e-13 K=2.62 tau=1.0685844340773973e-07 off=-0.1

*Grain_238:
XU_238 in out fe_tanh Vc=0.8227241003637082 Qo=7.074306885472911e-13 K=2.62 tau=9.53723156760807e-08 off=-0.1

*Grain_239:
XU_239 in out fe_tanh Vc=0.414349520251386 Qo=2.9002157243746187e-13 K=2.62 tau=7.97043057986304e-08 off=-0.1

*Grain_240:
XU_240 in out fe_tanh Vc=0.6543253964344135 Qo=5.25273293477712e-13 K=2.62 tau=8.479740110009681e-08 off=-0.1

*Grain_241:
XU_241 in out fe_tanh Vc=0.057356002941954365 Qo=2.218226821833358e-14 K=2.62 tau=7.457618354726614e-08 off=-0.1

*Grain_242:
XU_242 in out fe_tanh Vc=0.8876432222895947 Qo=7.808423937161502e-13 K=2.62 tau=1.1425744565075558e-07 off=-0.1

*Grain_243:
XU_243 in out fe_tanh Vc=0.41630350693125906 Qo=2.918008150627689e-13 K=2.62 tau=9.461496087987213e-08 off=-0.1

*Grain_244:
XU_244 in out fe_tanh Vc=0.6586580618350976 Qo=5.297993557601956e-13 K=2.62 tau=8.906912775272348e-08 off=-0.1

*Grain_245:
XU_245 in out fe_tanh Vc=0.43740240005473197 Qo=3.1117086036120676e-13 K=2.62 tau=1.0115201454695113e-07 off=-0.1

*Grain_246:
XU_246 in out fe_tanh Vc=0.435344220809468 Qo=3.092687429245935e-13 K=2.62 tau=1.0217839839919251e-07 off=-0.1

*Grain_247:
XU_247 in out fe_tanh Vc=0.3092116456136191 Qo=1.9823758809902345e-13 K=2.62 tau=9.742085193576366e-08 off=-0.1

*Grain_248:
XU_248 in out fe_tanh Vc=0.45837713436860494 Qo=3.3070688697638915e-13 K=2.62 tau=1.0504279576226138e-07 off=-0.1

*Grain_249:
XU_249 in out fe_tanh Vc=0.21767580788707835 Qo=1.256049123855874e-13 K=2.62 tau=1.0222744076537703e-07 off=-0.1

*Grain_250:
XU_250 in out fe_tanh Vc=0.4717580830956455 Qo=3.433116693296572e-13 K=2.62 tau=1.206091411163463e-07 off=-0.1

*Grain_251:
XU_251 in out fe_tanh Vc=0.6785484483104056 Qo=5.506916997141054e-13 K=2.62 tau=9.624545838509405e-08 off=-0.1

*Grain_252:
XU_252 in out fe_tanh Vc=0.2921838408568582 Qo=1.8416473069500212e-13 K=2.62 tau=7.567065432221147e-08 off=-0.1

*Grain_253:
XU_253 in out fe_tanh Vc=0.3813868105870212 Qo=2.603926858800039e-13 K=2.62 tau=1.0244732258759756e-07 off=-0.1

*Grain_254:
XU_254 in out fe_tanh Vc=0.44527647836803336 Qo=3.184726128034825e-13 K=2.62 tau=1.1321422153926605e-07 off=-0.1

*Grain_255:
XU_255 in out fe_tanh Vc=0.30039614538714576 Qo=1.9092204288593687e-13 K=2.62 tau=1.029900369438668e-07 off=-0.1

*Grain_256:
XU_256 in out fe_tanh Vc=0.45999687608876155 Qo=3.322268721817917e-13 K=2.62 tau=1.1575629648903273e-07 off=-0.1

*Grain_257:
XU_257 in out fe_tanh Vc=0.04424285556712926 Qo=1.5828855164179794e-14 K=2.62 tau=9.536650373229895e-08 off=-0.1

*Grain_258:
XU_258 in out fe_tanh Vc=0.20613859251307445 Qo=1.1702011182029688e-13 K=2.62 tau=1.1350332824218131e-07 off=-0.1

*Grain_259:
XU_259 in out fe_tanh Vc=0.5510960659283924 Qo=4.201930979307382e-13 K=2.62 tau=9.769396746511375e-08 off=-0.1

*Grain_260:
XU_260 in out fe_tanh Vc=0.1522374933332947 Qo=7.89099053085628e-14 K=2.62 tau=1.1206591412527204e-07 off=-0.1

*Grain_261:
XU_261 in out fe_tanh Vc=1.005535454381053 Qo=9.182691940891402e-13 K=2.62 tau=1.0213409986000806e-07 off=-0.1

*Grain_262:
XU_262 in out fe_tanh Vc=0.7061591784952755 Qo=5.799984077121173e-13 K=2.62 tau=8.385922445747282e-08 off=-0.1

*Grain_263:
XU_263 in out fe_tanh Vc=0.544969506665893 Qo=4.141305541347479e-13 K=2.62 tau=1.1527165101152963e-07 off=-0.1

*Grain_264:
XU_264 in out fe_tanh Vc=0.7162621389140291 Qo=5.908088664737112e-13 K=2.62 tau=9.610151223111283e-08 off=-0.1

*Grain_265:
XU_265 in out fe_tanh Vc=0.45655508834586556 Qo=3.2899898192413925e-13 K=2.62 tau=9.711472933664357e-08 off=-0.1

*Grain_266:
XU_266 in out fe_tanh Vc=0.5845545049395873 Qo=4.5365523390322663e-13 K=2.62 tau=8.58831972448947e-08 off=-0.1

*Grain_267:
XU_267 in out fe_tanh Vc=-0.25883821760679326 Qo=1.573223159840978e-13 K=2.62 tau=1.0111538693707894e-07 off=-0.1

*Grain_268:
XU_268 in out fe_tanh Vc=0.9163942540527894 Qo=8.138801849150683e-13 K=2.62 tau=1.0610598452630207e-07 off=-0.1

*Grain_269:
XU_269 in out fe_tanh Vc=0.2571617066089741 Qo=1.559989227753247e-13 K=2.62 tau=1.2605952846527953e-07 off=-0.1

*Grain_270:
XU_270 in out fe_tanh Vc=0.7047299545801826 Qo=5.784728245400323e-13 K=2.62 tau=1.0130058553133974e-07 off=-0.1

*Grain_271:
XU_271 in out fe_tanh Vc=0.5839434763073503 Qo=4.5303886926991306e-13 K=2.62 tau=1.0891617245270365e-07 off=-0.1

*Grain_272:
XU_272 in out fe_tanh Vc=-0.07321264276280726 Qo=3.046599170492992e-14 K=2.62 tau=7.957333503387856e-08 off=-0.1

*Grain_273:
XU_273 in out fe_tanh Vc=0.3126797267043835 Qo=2.011328702598105e-13 K=2.62 tau=1.0530406459510848e-07 off=-0.1

*Grain_274:
XU_274 in out fe_tanh Vc=0.19819983959530002 Qo=1.1119562460842909e-13 K=2.62 tau=9.433075966321516e-08 off=-0.1

*Grain_275:
XU_275 in out fe_tanh Vc=0.4223908251463657 Qo=2.973597818695393e-13 K=2.62 tau=1.1685758502526423e-07 off=-0.1

*Grain_276:
XU_276 in out fe_tanh Vc=0.341022388267083 Qo=2.2514959466623637e-13 K=2.62 tau=9.899621594761126e-08 off=-0.1

*Grain_277:
XU_277 in out fe_tanh Vc=0.5904303160415435 Qo=4.595922043384351e-13 K=2.62 tau=1.1185597353718108e-07 off=-0.1

*Grain_278:
XU_278 in out fe_tanh Vc=0.4358088100463545 Qo=3.09697869330821e-13 K=2.62 tau=1.0052373964608845e-07 off=-0.1

*Grain_279:
XU_279 in out fe_tanh Vc=0.536053522459615 Qo=4.0534424449415467e-13 K=2.62 tau=1.0706921947381991e-07 off=-0.1

*Grain_280:
XU_280 in out fe_tanh Vc=0.5363148317409933 Qo=4.056011336641524e-13 K=2.62 tau=9.161278084444955e-08 off=-0.1

*Grain_281:
XU_281 in out fe_tanh Vc=0.29460501959668384 Qo=1.8615109505881758e-13 K=2.62 tau=9.289937379823495e-08 off=-0.1

*Grain_282:
XU_282 in out fe_tanh Vc=0.5017961484532732 Qo=3.7199656620710394e-13 K=2.62 tau=9.82154864665418e-08 off=-0.1

*Grain_283:
XU_283 in out fe_tanh Vc=0.4773856708768908 Qo=3.486451301109624e-13 K=2.62 tau=8.153719938907052e-08 off=-0.1

*Grain_284:
XU_284 in out fe_tanh Vc=0.7125984160893754 Qo=5.8688325577656e-13 K=2.62 tau=1.0131032953311832e-07 off=-0.1

*Grain_285:
XU_285 in out fe_tanh Vc=0.11802567915567402 Qo=5.667909028127208e-14 K=2.62 tau=9.157379253454947e-08 off=-0.1

*Grain_286:
XU_286 in out fe_tanh Vc=0.1737218825154481 Qo=9.368375623785057e-14 K=2.62 tau=8.285137880904627e-08 off=-0.1

*Grain_287:
XU_287 in out fe_tanh Vc=0.2928495601001087 Qo=1.847104044342441e-13 K=2.62 tau=9.972127262817941e-08 off=-0.1

*Grain_288:
XU_288 in out fe_tanh Vc=0.23711568140659206 Qo=1.4037887897953123e-13 K=2.62 tau=1.1414001768211149e-07 off=-0.1

*Grain_289:
XU_289 in out fe_tanh Vc=-0.7337982337400476 Qo=6.096815758181864e-13 K=2.62 tau=9.228103665821182e-08 off=-0.1

*Grain_290:
XU_290 in out fe_tanh Vc=0.6084318400455884 Qo=4.778910791492442e-13 K=2.62 tau=1.1715683053469108e-07 off=-0.1

*Grain_291:
XU_291 in out fe_tanh Vc=0.13646987730697968 Qo=6.845438165617366e-14 K=2.62 tau=9.42916849290619e-08 off=-0.1

*Grain_292:
XU_292 in out fe_tanh Vc=0.2646108006741655 Qo=1.618986574637938e-13 K=2.62 tau=8.834148512908943e-08 off=-0.1

*Grain_293:
XU_293 in out fe_tanh Vc=0.45900297629245657 Qo=3.312939939045141e-13 K=2.62 tau=1.1449822109787829e-07 off=-0.1

*Grain_294:
XU_294 in out fe_tanh Vc=0.40832527603901086 Qo=2.8455194209982395e-13 K=2.62 tau=1.0487399712210033e-07 off=-0.1

*Grain_295:
XU_295 in out fe_tanh Vc=-0.006265552363578009 Qo=1.2470980021861863e-15 K=2.62 tau=9.3059832564423e-08 off=-0.1

*Grain_296:
XU_296 in out fe_tanh Vc=0.2113572687233761 Qo=1.2088592972714765e-13 K=2.62 tau=9.504637079581567e-08 off=-0.1

*Grain_297:
XU_297 in out fe_tanh Vc=0.3205833164016311 Qo=2.077670162713786e-13 K=2.62 tau=1.1261987096487511e-07 off=-0.1

*Grain_298:
XU_298 in out fe_tanh Vc=0.5841741287286741 Qo=4.5327151321418676e-13 K=2.62 tau=8.190960465544555e-08 off=-0.1

*Grain_299:
XU_299 in out fe_tanh Vc=0.5131313702623796 Qo=3.829574708439796e-13 K=2.62 tau=8.06110345997665e-08 off=-0.1

*Grain_300:
XU_300 in out fe_tanh Vc=1.2626653085456856 Qo=1.2346052899305152e-12 K=2.62 tau=1.124456144642874e-07 off=-0.1

*Grain_301:
XU_301 in out fe_tanh Vc=0.011853501937194255 Qo=2.8566306259116557e-15 K=2.62 tau=8.753546017455338e-08 off=-0.1

*Grain_302:
XU_302 in out fe_tanh Vc=0.2033244078030835 Qo=1.149475664598739e-13 K=2.62 tau=1.0408441920915759e-07 off=-0.1

*Grain_303:
XU_303 in out fe_tanh Vc=0.8123766597659549 Qo=6.958859672418413e-13 K=2.62 tau=9.096288130343175e-08 off=-0.1

*Grain_304:
XU_304 in out fe_tanh Vc=0.3679000828286175 Qo=2.4848619261006056e-13 K=2.62 tau=1.0579143474860815e-07 off=-0.1

*Grain_305:
XU_305 in out fe_tanh Vc=0.7508231540873548 Qo=6.281340908430464e-13 K=2.62 tau=9.441407541172287e-08 off=-0.1

*Grain_306:
XU_306 in out fe_tanh Vc=0.6468307291806248 Qo=5.174653180331251e-13 K=2.62 tau=9.72040793595012e-08 off=-0.1

*Grain_307:
XU_307 in out fe_tanh Vc=0.35530461307065947 Qo=2.3748408486336483e-13 K=2.62 tau=1.0579062387385838e-07 off=-0.1

*Grain_308:
XU_308 in out fe_tanh Vc=-0.16918265107403185 Qo=9.051404722260461e-14 K=2.62 tau=9.69498851591867e-08 off=-0.1

*Grain_309:
XU_309 in out fe_tanh Vc=0.34938431512794144 Qo=2.32352760255718e-13 K=2.62 tau=1.0074882710521643e-07 off=-0.1

*Grain_310:
XU_310 in out fe_tanh Vc=0.3682135972367159 Qo=2.4876150688647565e-13 K=2.62 tau=8.825437043315195e-08 off=-0.1

*Grain_311:
XU_311 in out fe_tanh Vc=0.43239430380181904 Qo=3.065472071349826e-13 K=2.62 tau=8.122624409572846e-08 off=-0.1

*Grain_312:
XU_312 in out fe_tanh Vc=0.26083107359935614 Qo=1.58898770966927e-13 K=2.62 tau=1.0122215256904532e-07 off=-0.1

*Grain_313:
XU_313 in out fe_tanh Vc=0.6943969077281416 Qo=5.67470803732527e-13 K=2.62 tau=1.0645235704413635e-07 off=-0.1

*Grain_314:
XU_314 in out fe_tanh Vc=0.21319594372632447 Qo=1.222548308829187e-13 K=2.62 tau=1.1032309512236314e-07 off=-0.1

*Grain_315:
XU_315 in out fe_tanh Vc=0.2375384432605354 Qo=1.4070433830760608e-13 K=2.62 tau=1.0934264592695712e-07 off=-0.1

*Grain_316:
XU_316 in out fe_tanh Vc=0.861819995710438 Qo=7.514411025686883e-13 K=2.62 tau=9.317735047142634e-08 off=-0.1

*Grain_317:
XU_317 in out fe_tanh Vc=0.3392937911010088 Qo=2.236670946648882e-13 K=2.62 tau=9.947567255643209e-08 off=-0.1

*Grain_318:
XU_318 in out fe_tanh Vc=0.1491422232972459 Qo=7.683059689795119e-14 K=2.62 tau=1.0580565516649288e-07 off=-0.1

*Grain_319:
XU_319 in out fe_tanh Vc=0.5723150816728892 Qo=4.4134596277575545e-13 K=2.62 tau=1.040467511329435e-07 off=-0.1

*Grain_320:
XU_320 in out fe_tanh Vc=0.8210880518867458 Qo=7.056024217471174e-13 K=2.62 tau=9.497533533253243e-08 off=-0.1

*Grain_321:
XU_321 in out fe_tanh Vc=0.2981081832626744 Qo=1.8903380563372255e-13 K=2.62 tau=9.585842946748612e-08 off=-0.1

*Grain_322:
XU_322 in out fe_tanh Vc=0.33577298463944005 Qo=2.2065454980020806e-13 K=2.62 tau=1.0233458891917066e-07 off=-0.1

*Grain_323:
XU_323 in out fe_tanh Vc=0.2436454960423581 Qo=1.4542508096135317e-13 K=2.62 tau=1.094019571001224e-07 off=-0.1

*Grain_324:
XU_324 in out fe_tanh Vc=0.26374937269619525 Qo=1.6121382282496971e-13 K=2.62 tau=1.0500836731885707e-07 off=-0.1

*Grain_325:
XU_325 in out fe_tanh Vc=0.11792064289007809 Qo=5.6613525442547144e-14 K=2.62 tau=9.634753104970657e-08 off=-0.1

*Grain_326:
XU_326 in out fe_tanh Vc=0.11785845143552776 Qo=5.657471308121776e-14 K=2.62 tau=8.825120273586315e-08 off=-0.1

*Grain_327:
XU_327 in out fe_tanh Vc=0.7637367053408826 Qo=6.42214597502429e-13 K=2.62 tau=1.042211372586319e-07 off=-0.1

*Grain_328:
XU_328 in out fe_tanh Vc=0.2945004115968982 Qo=1.860651718337544e-13 K=2.62 tau=1.0806474862378597e-07 off=-0.1

*Grain_329:
XU_329 in out fe_tanh Vc=0.33830976752546055 Qo=2.2282417547916082e-13 K=2.62 tau=9.422865620949406e-08 off=-0.1

*Grain_330:
XU_330 in out fe_tanh Vc=0.5130342152359268 Qo=3.828632128328141e-13 K=2.62 tau=1.0594139411746478e-07 off=-0.1

*Grain_331:
XU_331 in out fe_tanh Vc=0.297676794789093 Qo=1.8867826998119725e-13 K=2.62 tau=8.346214721733165e-08 off=-0.1

*Grain_332:
XU_332 in out fe_tanh Vc=0.5736738805987209 Qo=4.427086527728091e-13 K=2.62 tau=8.816612932373423e-08 off=-0.1

*Grain_333:
XU_333 in out fe_tanh Vc=0.21303309963016187 Qo=1.221334493293748e-13 K=2.62 tau=1.0959065266117243e-07 off=-0.1

*Grain_334:
XU_334 in out fe_tanh Vc=0.3630556759687523 Qo=2.4424102311887205e-13 K=2.62 tau=9.349952524107199e-08 off=-0.1

*Grain_335:
XU_335 in out fe_tanh Vc=0.3226745311957573 Qo=2.0953062310913472e-13 K=2.62 tau=8.609055188765838e-08 off=-0.1

*Grain_336:
XU_336 in out fe_tanh Vc=0.29832531909155563 Qo=1.8921281999034935e-13 K=2.62 tau=9.931335897868233e-08 off=-0.1

*Grain_337:
XU_337 in out fe_tanh Vc=-0.18031501503053515 Qo=9.833199956627555e-14 K=2.62 tau=1.098428185814212e-07 off=-0.1

*Grain_338:
XU_338 in out fe_tanh Vc=0.19206559824386277 Qo=1.0674262255720927e-13 K=2.62 tau=1.1442711746340754e-07 off=-0.1

*Grain_339:
XU_339 in out fe_tanh Vc=0.1300331985441453 Qo=6.428711396634762e-14 K=2.62 tau=1.0220771179378604e-07 off=-0.1

*Grain_340:
XU_340 in out fe_tanh Vc=0.21102677872165423 Qo=1.2064025621625877e-13 K=2.62 tau=8.772464876828037e-08 off=-0.1

*Grain_341:
XU_341 in out fe_tanh Vc=-0.016062383310824213 Qo=4.240395761839111e-15 K=2.62 tau=1.231550823243597e-07 off=-0.1

*Grain_342:
XU_342 in out fe_tanh Vc=0.49711803759334783 Qo=3.6749445317681125e-13 K=2.62 tau=9.7870299968881e-08 off=-0.1

*Grain_343:
XU_343 in out fe_tanh Vc=0.34277689224611846 Qo=2.2665662020906649e-13 K=2.62 tau=9.905846782687016e-08 off=-0.1

*Grain_344:
XU_344 in out fe_tanh Vc=0.2288536608035089 Qo=1.3405364694524864e-13 K=2.62 tau=1.0102875062524803e-07 off=-0.1

*Grain_345:
XU_345 in out fe_tanh Vc=0.004821949341254517 Qo=8.872435419272148e-16 K=2.62 tau=1.1810516911398246e-07 off=-0.1

*Grain_346:
XU_346 in out fe_tanh Vc=-0.013928504968468813 Qo=3.5231348381736734e-15 K=2.62 tau=1.0342361630806785e-07 off=-0.1

*Grain_347:
XU_347 in out fe_tanh Vc=0.5485375288030069 Qo=4.1765882254954765e-13 K=2.62 tau=1.1144225680890813e-07 off=-0.1

*Grain_348:
XU_348 in out fe_tanh Vc=0.22219882866845836 Qo=1.2900831569105438e-13 K=2.62 tau=1.0500311228239486e-07 off=-0.1

*Grain_349:
XU_349 in out fe_tanh Vc=0.12463555334032689 Qo=6.083982279403575e-14 K=2.62 tau=1.0053618137835756e-07 off=-0.1

*Grain_350:
XU_350 in out fe_tanh Vc=0.04788145339278671 Qo=1.7541669823626374e-14 K=2.62 tau=9.004089864471696e-08 off=-0.1

*Grain_351:
XU_351 in out fe_tanh Vc=0.24719958849889517 Qo=1.4818883265902895e-13 K=2.62 tau=9.769625389595382e-08 off=-0.1

*Grain_352:
XU_352 in out fe_tanh Vc=0.5494344337752656 Qo=4.1854681967646793e-13 K=2.62 tau=9.502533333165736e-08 off=-0.1

*Grain_353:
XU_353 in out fe_tanh Vc=0.7582462105830593 Qo=6.362191448068945e-13 K=2.62 tau=1.0618309893601426e-07 off=-0.1

*Grain_354:
XU_354 in out fe_tanh Vc=0.34079857566347427 Qo=2.2495751853179288e-13 K=2.62 tau=1.0742326607958406e-07 off=-0.1

*Grain_355:
XU_355 in out fe_tanh Vc=0.08728892863904775 Qo=3.829131864450153e-14 K=2.62 tau=8.040095847343754e-08 off=-0.1

*Grain_356:
XU_356 in out fe_tanh Vc=0.7206612801239431 Qo=5.955304275429012e-13 K=2.62 tau=1.0068201512602842e-07 off=-0.1

*Grain_357:
XU_357 in out fe_tanh Vc=0.4213435147603791 Qo=2.964016509209108e-13 K=2.62 tau=1.152102768272791e-07 off=-0.1

*Grain_358:
XU_358 in out fe_tanh Vc=0.06772539050064486 Qo=2.753153232348076e-14 K=2.62 tau=9.617211034146124e-08 off=-0.1

*Grain_359:
XU_359 in out fe_tanh Vc=0.26967213033111925 Qo=1.659358774520404e-13 K=2.62 tau=7.775531696335146e-08 off=-0.1

*Grain_360:
XU_360 in out fe_tanh Vc=0.7140904086505419 Qo=5.884811689717369e-13 K=2.62 tau=9.306153447619829e-08 off=-0.1

*Grain_361:
XU_361 in out fe_tanh Vc=0.42636148630388776 Qo=3.0099880276914456e-13 K=2.62 tau=8.859929288314671e-08 off=-0.1

*Grain_362:
XU_362 in out fe_tanh Vc=0.4577596751522354 Qo=3.301278795494606e-13 K=2.62 tau=9.877984440457856e-08 off=-0.1

*Grain_363:
XU_363 in out fe_tanh Vc=0.11163151810550082 Qo=5.272010791391258e-14 K=2.62 tau=1.2762655953820264e-07 off=-0.1

*Grain_364:
XU_364 in out fe_tanh Vc=0.055565835619945825 Qo=2.1286468439287843e-14 K=2.62 tau=8.967696781478957e-08 off=-0.1

*Grain_365:
XU_365 in out fe_tanh Vc=0.5095237415909468 Qo=3.794610140761776e-13 K=2.62 tau=8.50145454715572e-08 off=-0.1

*Grain_366:
XU_366 in out fe_tanh Vc=0.24829629704133457 Qo=1.4904407842263732e-13 K=2.62 tau=9.277864404493813e-08 off=-0.1

*Grain_367:
XU_367 in out fe_tanh Vc=0.8989074967038149 Qo=7.937484925554257e-13 K=2.62 tau=9.634968961234223e-08 off=-0.1

*Grain_368:
XU_368 in out fe_tanh Vc=-0.10148173431889473 Qo=4.6575513884983817e-14 K=2.62 tau=1.1269951966150654e-07 off=-0.1

*Grain_369:
XU_369 in out fe_tanh Vc=-0.4198320170177736 Qo=2.95020118098658e-13 K=2.62 tau=9.072306849224374e-08 off=-0.1

*Grain_370:
XU_370 in out fe_tanh Vc=0.5833360179988606 Qo=4.524262979025159e-13 K=2.62 tau=8.76911352818578e-08 off=-0.1

*Grain_371:
XU_371 in out fe_tanh Vc=0.7886852894836982 Qo=6.696197787198488e-13 K=2.62 tau=1.0287151703383451e-07 off=-0.1

*Grain_372:
XU_372 in out fe_tanh Vc=-0.17135798410549308 Qo=9.202992288646571e-14 K=2.62 tau=9.858617329020096e-08 off=-0.1

*Grain_373:
XU_373 in out fe_tanh Vc=0.5317271794634801 Qo=4.01096551868813e-13 K=2.62 tau=1.0184793162976474e-07 off=-0.1

*Grain_374:
XU_374 in out fe_tanh Vc=0.5319784805984472 Qo=4.0134300177335144e-13 K=2.62 tau=1.215438985090348e-07 off=-0.1

*Grain_375:
XU_375 in out fe_tanh Vc=0.32902005121153477 Qo=2.1490300373729633e-13 K=2.62 tau=1.0303091937685117e-07 off=-0.1

*Grain_376:
XU_376 in out fe_tanh Vc=0.08640823183557444 Qo=3.7789840963380174e-14 K=2.62 tau=9.460529656779478e-08 off=-0.1

*Grain_377:
XU_377 in out fe_tanh Vc=0.275391908273711 Qo=1.7052573828502189e-13 K=2.62 tau=9.510670362092833e-08 off=-0.1

*Grain_378:
XU_378 in out fe_tanh Vc=0.430928439929473 Qo=3.051968976562779e-13 K=2.62 tau=1.0922524807291208e-07 off=-0.1

*Grain_379:
XU_379 in out fe_tanh Vc=0.13581189655819842 Qo=6.802562938473083e-14 K=2.62 tau=9.486712656090092e-08 off=-0.1

*Grain_380:
XU_380 in out fe_tanh Vc=0.013745161688249241 Qo=3.4629659335046257e-15 K=2.62 tau=9.40997303493926e-08 off=-0.1

*Grain_381:
XU_381 in out fe_tanh Vc=0.7670158994785071 Qo=6.458015557816627e-13 K=2.62 tau=1.0494153860504002e-07 off=-0.1

*Grain_382:
XU_382 in out fe_tanh Vc=0.7023124066314108 Qo=5.758943967846786e-13 K=2.62 tau=9.877372412884913e-08 off=-0.1

*Grain_383:
XU_383 in out fe_tanh Vc=0.37089841938229734 Qo=2.5112207297500545e-13 K=2.62 tau=1.0911660603587432e-07 off=-0.1

*Grain_384:
XU_384 in out fe_tanh Vc=0.12311134105429727 Qo=5.987436095516901e-14 K=2.62 tau=1.1302515241124444e-07 off=-0.1

*Grain_385:
XU_385 in out fe_tanh Vc=0.22325864802729836 Qo=1.29808815812136e-13 K=2.62 tau=9.617976619297404e-08 off=-0.1

*Grain_386:
XU_386 in out fe_tanh Vc=0.6820946870444147 Qo=5.544360709501366e-13 K=2.62 tau=9.422989195672418e-08 off=-0.1

*Grain_387:
XU_387 in out fe_tanh Vc=0.3535630315327012 Qo=2.359719134257965e-13 K=2.62 tau=1.0071202380034906e-07 off=-0.1

*Grain_388:
XU_388 in out fe_tanh Vc=-0.07515464563231128 Qo=3.1520709989140086e-14 K=2.62 tau=1.1281245333609462e-07 off=-0.1

*Grain_389:
XU_389 in out fe_tanh Vc=0.7053299783631131 Qo=5.791131894083632e-13 K=2.62 tau=1.0691370123218877e-07 off=-0.1

*Grain_390:
XU_390 in out fe_tanh Vc=0.25491411977010014 Qo=1.5422879656023435e-13 K=2.62 tau=8.783236655935502e-08 off=-0.1

*Grain_391:
XU_391 in out fe_tanh Vc=0.6177335183283267 Qo=4.874105523693875e-13 K=2.62 tau=9.960660194678804e-08 off=-0.1

*Grain_392:
XU_392 in out fe_tanh Vc=0.41575719617907386 Qo=2.913031077646381e-13 K=2.62 tau=1.0565716374188025e-07 off=-0.1

*Grain_393:
XU_393 in out fe_tanh Vc=-0.20954354497450467 Qo=1.19539100441834e-13 K=2.62 tau=8.929679214334954e-08 off=-0.1

*Grain_394:
XU_394 in out fe_tanh Vc=0.6757911406405384 Qo=5.477843906519823e-13 K=2.62 tau=9.306502424192202e-08 off=-0.1

*Grain_395:
XU_395 in out fe_tanh Vc=0.5842510926300506 Qo=4.5334914777764135e-13 K=2.62 tau=9.42659452909925e-08 off=-0.1

*Grain_396:
XU_396 in out fe_tanh Vc=0.3983032240215573 Qo=2.75506201307924e-13 K=2.62 tau=9.931695137828825e-08 off=-0.1

*Grain_397:
XU_397 in out fe_tanh Vc=0.74753403406893 Qo=6.245592886271952e-13 K=2.62 tau=9.080630889677631e-08 off=-0.1

*Grain_398:
XU_398 in out fe_tanh Vc=-0.052579833208292404 Qo=1.9811546393490492e-14 K=2.62 tau=1.1211809188700414e-07 off=-0.1

*Grain_399:
XU_399 in out fe_tanh Vc=-0.08115538502381436 Qo=3.4831000997064565e-14 K=2.62 tau=1.1175206015047127e-07 off=-0.1

*Grain_400:
XU_400 in out fe_tanh Vc=0.8793880775322327 Qo=7.714151355987777e-13 K=2.62 tau=9.653517281426361e-08 off=-0.1

*Grain_401:
XU_401 in out fe_tanh Vc=0.5158713100737204 Qo=3.8561791183582767e-13 K=2.62 tau=1.0433251944973498e-07 off=-0.1

*Grain_402:
XU_402 in out fe_tanh Vc=0.44237667600987257 Qo=3.157790383109858e-13 K=2.62 tau=1.005736204067935e-07 off=-0.1

*Grain_403:
XU_403 in out fe_tanh Vc=-0.05683908960795497 Qo=2.1922731134873392e-14 K=2.62 tau=9.353810645297551e-08 off=-0.1

*Grain_404:
XU_404 in out fe_tanh Vc=-0.05858089380148834 Qo=2.280007114680795e-14 K=2.62 tau=1.1186295752970992e-07 off=-0.1

*Grain_405:
XU_405 in out fe_tanh Vc=0.017613541296535473 Qo=4.780288379449755e-15 K=2.62 tau=1.0507287763081764e-07 off=-0.1

*Grain_406:
XU_406 in out fe_tanh Vc=0.49901812407362 Qo=3.6932152949453873e-13 K=2.62 tau=9.683598745972733e-08 off=-0.1

*Grain_407:
XU_407 in out fe_tanh Vc=0.18855894981876817 Qo=1.0421607348349068e-13 K=2.62 tau=9.771728354368239e-08 off=-0.1

*Grain_408:
XU_408 in out fe_tanh Vc=-0.11384345227358905 Qo=5.408214207431395e-14 K=2.62 tau=1.201773408085423e-07 off=-0.1

*Grain_409:
XU_409 in out fe_tanh Vc=0.12365842922291481 Qo=6.022048566060264e-14 K=2.62 tau=9.227378856429611e-08 off=-0.1

*Grain_410:
XU_410 in out fe_tanh Vc=0.2147166549477259 Qo=1.2338968710910512e-13 K=2.62 tau=8.504528836477671e-08 off=-0.1

*Grain_411:
XU_411 in out fe_tanh Vc=0.09708433788565929 Qo=4.396907562665817e-14 K=2.62 tau=8.606240221161385e-08 off=-0.1

*Grain_412:
XU_412 in out fe_tanh Vc=0.3004240289827964 Qo=1.9094508168793733e-13 K=2.62 tau=9.781796641693576e-08 off=-0.1

*Grain_413:
XU_413 in out fe_tanh Vc=0.711750139134945 Qo=5.859752046304074e-13 K=2.62 tau=1.1120583636692809e-07 off=-0.1

*Grain_414:
XU_414 in out fe_tanh Vc=0.7111243971660874 Qo=5.853055775207568e-13 K=2.62 tau=1.0340356580617822e-07 off=-0.1

*Grain_415:
XU_415 in out fe_tanh Vc=0.46675765473646097 Qo=3.3858857075232154e-13 K=2.62 tau=1.0825329786439526e-07 off=-0.1

*Grain_416:
XU_416 in out fe_tanh Vc=0.0532159950242968 Qo=2.012371942037936e-14 K=2.62 tau=1.1011863193083913e-07 off=-0.1

*Grain_417:
XU_417 in out fe_tanh Vc=0.9073440019682258 Qo=8.034465215993042e-13 K=2.62 tau=1.0780433965827969e-07 off=-0.1

*Grain_418:
XU_418 in out fe_tanh Vc=0.2641712787265318 Qo=1.615491541172029e-13 K=2.62 tau=9.999720155789516e-08 off=-0.1

*Grain_419:
XU_419 in out fe_tanh Vc=0.5519684938846164 Qo=4.2105806108486176e-13 K=2.62 tau=9.586355593670956e-08 off=-0.1

*Grain_420:
XU_420 in out fe_tanh Vc=-0.07176006501713816 Qo=2.968254131792472e-14 K=2.62 tau=1.0768499480481363e-07 off=-0.1

*Grain_421:
XU_421 in out fe_tanh Vc=0.4307683437050056 Qo=3.0504950522076246e-13 K=2.62 tau=1.0768420259518851e-07 off=-0.1

*Grain_422:
XU_422 in out fe_tanh Vc=0.6047143655397779 Qo=4.740987190950316e-13 K=2.62 tau=1.0001267437278997e-07 off=-0.1

*Grain_423:
XU_423 in out fe_tanh Vc=0.39443948584583277 Qo=2.7203695792169585e-13 K=2.62 tau=1.0782692602280641e-07 off=-0.1

*Grain_424:
XU_424 in out fe_tanh Vc=0.2013838011020936 Qo=1.135233777281735e-13 K=2.62 tau=8.521104414702302e-08 off=-0.1

*Grain_425:
XU_425 in out fe_tanh Vc=0.41313728207886685 Qo=2.8891900792578394e-13 K=2.62 tau=9.96838350392689e-08 off=-0.1

*Grain_426:
XU_426 in out fe_tanh Vc=0.4251007661804424 Qo=2.9984227507837467e-13 K=2.62 tau=1.1640305969277196e-07 off=-0.1

*Grain_427:
XU_427 in out fe_tanh Vc=0.5407314838468595 Qo=4.0994874801903523e-13 K=2.62 tau=9.093421602819482e-08 off=-0.1

*Grain_428:
XU_428 in out fe_tanh Vc=0.8735866364461402 Qo=7.648058247303831e-13 K=2.62 tau=9.528293419106082e-08 off=-0.1

*Grain_429:
XU_429 in out fe_tanh Vc=0.3210258785146768 Qo=2.0813995987468554e-13 K=2.62 tau=1.0803039811120323e-07 off=-0.1

*Grain_430:
XU_430 in out fe_tanh Vc=0.10797568415882652 Qo=5.0486720901497424e-14 K=2.62 tau=9.682663089375931e-08 off=-0.1

*Grain_431:
XU_431 in out fe_tanh Vc=0.09968098178465706 Qo=4.550398266807734e-14 K=2.62 tau=9.928302600548162e-08 off=-0.1

*Grain_432:
XU_432 in out fe_tanh Vc=0.7724461958837245 Qo=6.517516221580608e-13 K=2.62 tau=8.234859551570866e-08 off=-0.1

*Grain_433:
XU_433 in out fe_tanh Vc=0.38645217225518985 Qo=2.648975179827784e-13 K=2.62 tau=1.1790590740763608e-07 off=-0.1

*Grain_434:
XU_434 in out fe_tanh Vc=0.7730151527142939 Qo=6.523757657587278e-13 K=2.62 tau=1.0060853990045727e-07 off=-0.1

*Grain_435:
XU_435 in out fe_tanh Vc=-0.10060127344061165 Qo=4.6050879829709445e-14 K=2.62 tau=1.1618053888013434e-07 off=-0.1

*Grain_436:
XU_436 in out fe_tanh Vc=0.6401645241993845 Qo=5.105431983561727e-13 K=2.62 tau=1.0009230725898993e-07 off=-0.1

*Grain_437:
XU_437 in out fe_tanh Vc=0.28676640085330984 Qo=1.7973810383117722e-13 K=2.62 tau=8.688517234543842e-08 off=-0.1

*Grain_438:
XU_438 in out fe_tanh Vc=0.4978705186049695 Qo=3.6821777026669113e-13 K=2.62 tau=1.0790080299617516e-07 off=-0.1

*Grain_439:
XU_439 in out fe_tanh Vc=1.3243639019100355 Qo=1.3135994125397772e-12 K=2.62 tau=1.129310661984799e-07 off=-0.1

*Grain_440:
XU_440 in out fe_tanh Vc=0.2533160506326027 Qo=1.5297305198437223e-13 K=2.62 tau=1.0109167789783488e-07 off=-0.1

*Grain_441:
XU_441 in out fe_tanh Vc=-0.58831793794504 Qo=4.574557889891049e-13 K=2.62 tau=1.213411785972738e-07 off=-0.1

*Grain_442:
XU_442 in out fe_tanh Vc=0.3262972255003322 Qo=2.12593903266176e-13 K=2.62 tau=9.515257346953538e-08 off=-0.1

*Grain_443:
XU_443 in out fe_tanh Vc=0.19653071823792123 Qo=1.0997981483278151e-13 K=2.62 tau=8.589208031929749e-08 off=-0.1

*Grain_444:
XU_444 in out fe_tanh Vc=0.4422429880933071 Qo=3.1565498541833393e-13 K=2.62 tau=1.1013130238785858e-07 off=-0.1

*Grain_445:
XU_445 in out fe_tanh Vc=0.6065594847022913 Qo=4.759801351704962e-13 K=2.62 tau=9.262948247633973e-08 off=-0.1

*Grain_446:
XU_446 in out fe_tanh Vc=0.27275499628516686 Qo=1.6840614694346137e-13 K=2.62 tau=1.011795798797566e-07 off=-0.1

*Grain_447:
XU_447 in out fe_tanh Vc=1.4520706750228487 Qo=1.4805991362447703e-12 K=2.62 tau=1.0934439369070055e-07 off=-0.1

*Grain_448:
XU_448 in out fe_tanh Vc=0.9450972591412089 Qo=8.471744808947238e-13 K=2.62 tau=1.071048780016799e-07 off=-0.1

*Grain_449:
XU_449 in out fe_tanh Vc=-0.12738705937648265 Qo=6.259163793215766e-14 K=2.62 tau=7.572970357428585e-08 off=-0.1

*Grain_450:
XU_450 in out fe_tanh Vc=0.7203016682987387 Qo=5.95144133890746e-13 K=2.62 tau=9.827032506900543e-08 off=-0.1

*Grain_451:
XU_451 in out fe_tanh Vc=0.06171991947503447 Qo=2.440092929139887e-14 K=2.62 tau=8.77990274677669e-08 off=-0.1

*Grain_452:
XU_452 in out fe_tanh Vc=0.7279006914407693 Qo=6.033192492153077e-13 K=2.62 tau=1.0530580261169973e-07 off=-0.1

*Grain_453:
XU_453 in out fe_tanh Vc=0.21754917466884938 Qo=1.2550992858308072e-13 K=2.62 tau=8.288389864038382e-08 off=-0.1

*Grain_454:
XU_454 in out fe_tanh Vc=0.2822801798979247 Qo=1.7609130485367647e-13 K=2.62 tau=9.304435058074894e-08 off=-0.1

*Grain_455:
XU_455 in out fe_tanh Vc=0.2665627248954364 Qo=1.634529094760846e-13 K=2.62 tau=8.96822219263284e-08 off=-0.1

*Grain_456:
XU_456 in out fe_tanh Vc=0.5383446287909271 Qo=4.0759787397943763e-13 K=2.62 tau=1.0469061761842309e-07 off=-0.1

*Grain_457:
XU_457 in out fe_tanh Vc=0.5135045853165247 Qo=3.8331960697421485e-13 K=2.62 tau=1.006186395588083e-07 off=-0.1

*Grain_458:
XU_458 in out fe_tanh Vc=0.9357483668964758 Qo=8.362963698438379e-13 K=2.62 tau=1.0021206241753275e-07 off=-0.1

*Grain_459:
XU_459 in out fe_tanh Vc=0.13193096142573896 Qo=6.550948057509549e-14 K=2.62 tau=9.505005669013593e-08 off=-0.1

*Grain_460:
XU_460 in out fe_tanh Vc=0.17403415612519052 Qo=9.390273673597336e-14 K=2.62 tau=9.99333717466439e-08 off=-0.1

*Grain_461:
XU_461 in out fe_tanh Vc=0.8330679590433455 Qo=7.190150336791945e-13 K=2.62 tau=9.254707440950552e-08 off=-0.1

*Grain_462:
XU_462 in out fe_tanh Vc=0.7649329072657305 Qo=6.435225330441951e-13 K=2.62 tau=1.0364702521882891e-07 off=-0.1

*Grain_463:
XU_463 in out fe_tanh Vc=0.30178777230348686 Qo=1.920726558125531e-13 K=2.62 tau=9.502090385670933e-08 off=-0.1

*Grain_464:
XU_464 in out fe_tanh Vc=0.37761797609996905 Qo=2.570525217410584e-13 K=2.62 tau=9.877058923502285e-08 off=-0.1

*Grain_465:
XU_465 in out fe_tanh Vc=0.6747252162537909 Qo=5.466614311159646e-13 K=2.62 tau=9.362960939973786e-08 off=-0.1

*Grain_466:
XU_466 in out fe_tanh Vc=0.21275326865212874 Qo=1.2192493251862109e-13 K=2.62 tau=1.0402994040464956e-07 off=-0.1

*Grain_467:
XU_467 in out fe_tanh Vc=0.47143758813213293 Qo=3.430084970348628e-13 K=2.62 tau=1.2179088488092304e-07 off=-0.1

*Grain_468:
XU_468 in out fe_tanh Vc=0.8429124604678154 Qo=7.300802943134778e-13 K=2.62 tau=9.466627759701293e-08 off=-0.1

*Grain_469:
XU_469 in out fe_tanh Vc=0.5324998617526202 Qo=4.018544293459633e-13 K=2.62 tau=9.95121161380363e-08 off=-0.1

*Grain_470:
XU_470 in out fe_tanh Vc=0.3364068933531768 Qo=2.2119625140778834e-13 K=2.62 tau=1.0809717667265387e-07 off=-0.1

*Grain_471:
XU_471 in out fe_tanh Vc=0.8576335375648719 Qo=7.466992116344994e-13 K=2.62 tau=8.816282395510814e-08 off=-0.1

*Grain_472:
XU_472 in out fe_tanh Vc=0.30152435751960277 Qo=1.9185473910737737e-13 K=2.62 tau=1.1775127192681062e-07 off=-0.1

*Grain_473:
XU_473 in out fe_tanh Vc=0.7053833941338713 Qo=5.79170204378128e-13 K=2.62 tau=9.665406556614847e-08 off=-0.1

*Grain_474:
XU_474 in out fe_tanh Vc=0.6642302207775606 Qo=5.356333761305668e-13 K=2.62 tau=9.832852222495569e-08 off=-0.1

*Grain_475:
XU_475 in out fe_tanh Vc=0.49263248433198215 Qo=3.6318957177258116e-13 K=2.62 tau=1.1669000334772024e-07 off=-0.1

*Grain_476:
XU_476 in out fe_tanh Vc=-0.03918258108792699 Qo=1.3516814812664418e-14 K=2.62 tau=8.857630693551803e-08 off=-0.1

*Grain_477:
XU_477 in out fe_tanh Vc=-0.08625978247423921 Qo=3.7705462880313664e-14 K=2.62 tau=9.187378363229146e-08 off=-0.1

*Grain_478:
XU_478 in out fe_tanh Vc=0.4442670836337011 Qo=3.175344052058354e-13 K=2.62 tau=9.847260466795036e-08 off=-0.1

*Grain_479:
XU_479 in out fe_tanh Vc=0.26393609846625105 Qo=1.6136221280019898e-13 K=2.62 tau=1.1247895843086405e-07 off=-0.1

*Grain_480:
XU_480 in out fe_tanh Vc=1.3072730066851888 Qo=1.2916046273262366e-12 K=2.62 tau=1.0530105353351754e-07 off=-0.1

*Grain_481:
XU_481 in out fe_tanh Vc=0.6419605197684203 Qo=5.124060235807981e-13 K=2.62 tau=1.0186706067821274e-07 off=-0.1

*Grain_482:
XU_482 in out fe_tanh Vc=0.31471800639437547 Qo=2.0283900868530535e-13 K=2.62 tau=8.423522520447147e-08 off=-0.1

*Grain_483:
XU_483 in out fe_tanh Vc=0.6973203033601411 Qo=5.70578514482884e-13 K=2.62 tau=8.900022497327571e-08 off=-0.1

*Grain_484:
XU_484 in out fe_tanh Vc=0.28562490057641504 Qo=1.788085562345557e-13 K=2.62 tau=1.0002667558143294e-07 off=-0.1

*Grain_485:
XU_485 in out fe_tanh Vc=0.5725729984023294 Qo=4.41604543523159e-13 K=2.62 tau=1.1613338989302833e-07 off=-0.1

*Grain_486:
XU_486 in out fe_tanh Vc=0.2562225782240928 Qo=1.5525872896098143e-13 K=2.62 tau=1.2517996512173207e-07 off=-0.1

*Grain_487:
XU_487 in out fe_tanh Vc=0.47420864543916474 Qo=3.456318199324328e-13 K=2.62 tau=1.0301507505349199e-07 off=-0.1

*Grain_488:
XU_488 in out fe_tanh Vc=0.6676615000225894 Qo=5.392332261097561e-13 K=2.62 tau=9.696843774239123e-08 off=-0.1

*Grain_489:
XU_489 in out fe_tanh Vc=0.7726186236572243 Qo=6.519407602464709e-13 K=2.62 tau=1.0321369931049511e-07 off=-0.1

*Grain_490:
XU_490 in out fe_tanh Vc=0.506244737899774 Qo=3.762894905975575e-13 K=2.62 tau=1.0319412517375667e-07 off=-0.1

*Grain_491:
XU_491 in out fe_tanh Vc=1.1726552284341576 Qo=1.1214369409278627e-12 K=2.62 tau=9.041505938196512e-08 off=-0.1

*Grain_492:
XU_492 in out fe_tanh Vc=0.37631485711109053 Qo=2.5589994038822633e-13 K=2.62 tau=1.1413241134693268e-07 off=-0.1

*Grain_493:
XU_493 in out fe_tanh Vc=1.0965836062841818 Qo=1.027797800846485e-12 K=2.62 tau=8.960849497679768e-08 off=-0.1

*Grain_494:
XU_494 in out fe_tanh Vc=0.5483673146363368 Qo=4.174903480585851e-13 K=2.62 tau=1.0914655462038751e-07 off=-0.1

*Grain_495:
XU_495 in out fe_tanh Vc=0.04794398202711403 Qo=1.7571455738324587e-14 K=2.62 tau=1.0550735850247751e-07 off=-0.1

*Grain_496:
XU_496 in out fe_tanh Vc=0.44331501016904457 Qo=3.166500621554823e-13 K=2.62 tau=1.049086527491687e-07 off=-0.1

*Grain_497:
XU_497 in out fe_tanh Vc=-0.054951851983115474 Qo=2.0981205818324712e-14 K=2.62 tau=1.072261508758823e-07 off=-0.1

*Grain_498:
XU_498 in out fe_tanh Vc=0.771706393422595 Qo=6.509402677565191e-13 K=2.62 tau=1.0096846728996531e-07 off=-0.1

*Grain_499:
XU_499 in out fe_tanh Vc=0.30365435792852435 Qo=1.9361847013910677e-13 K=2.62 tau=1.000436292895731e-07 off=-0.1

*Grain_500:
XU_500 in out fe_tanh Vc=0.6003082213819882 Qo=4.696128683540007e-13 K=2.62 tau=1.0132212017893536e-07 off=-0.1

*Grain_501:
XU_501 in out fe_tanh Vc=0.6329495820075207 Qo=5.030756106739933e-13 K=2.62 tau=9.659862028772886e-08 off=-0.1

*Grain_502:
XU_502 in out fe_tanh Vc=0.6651503522728699 Qo=5.365981653713293e-13 K=2.62 tau=9.891157168725487e-08 off=-0.1

*Grain_503:
XU_503 in out fe_tanh Vc=0.2873688806075546 Qo=1.8022916373616526e-13 K=2.62 tau=9.960203705372153e-08 off=-0.1

*Grain_504:
XU_504 in out fe_tanh Vc=0.6452367069123883 Qo=5.158081456796728e-13 K=2.62 tau=1.0364542062007308e-07 off=-0.1

*Grain_505:
XU_505 in out fe_tanh Vc=0.7048444875368791 Qo=5.785950452047076e-13 K=2.62 tau=1.2468584084518288e-07 off=-0.1

*Grain_506:
XU_506 in out fe_tanh Vc=0.4120950911378872 Qo=2.87971881594657e-13 K=2.62 tau=9.476560021336926e-08 off=-0.1

*Grain_507:
XU_507 in out fe_tanh Vc=0.36072113398753003 Qo=2.422013024663966e-13 K=2.62 tau=1.0847739468177522e-07 off=-0.1

*Grain_508:
XU_508 in out fe_tanh Vc=0.9202827091196346 Qo=8.183725455640728e-13 K=2.62 tau=1.0096406766438322e-07 off=-0.1

*Grain_509:
XU_509 in out fe_tanh Vc=0.39251153807430245 Qo=2.7030966000646585e-13 K=2.62 tau=1.0150848373305503e-07 off=-0.1

*Grain_510:
XU_510 in out fe_tanh Vc=0.11784543089539185 Qo=5.656658801731429e-14 K=2.62 tau=1.1150385473938189e-07 off=-0.1

*Grain_511:
XU_511 in out fe_tanh Vc=1.0390608824633136 Qo=9.582673788772983e-13 K=2.62 tau=8.627087103407276e-08 off=-0.1

*Grain_512:
XU_512 in out fe_tanh Vc=0.19451036052200577 Qo=1.085123005270662e-13 K=2.62 tau=1.0677457487852168e-07 off=-0.1

*Grain_513:
XU_513 in out fe_tanh Vc=0.056870044090408134 Qo=2.1938253214798454e-14 K=2.62 tau=8.375151141515546e-08 off=-0.1

*Grain_514:
XU_514 in out fe_tanh Vc=0.070006843668378 Qo=2.874326223635705e-14 K=2.62 tau=1.0019325872079855e-07 off=-0.1

*Grain_515:
XU_515 in out fe_tanh Vc=0.070321857963202 Qo=2.891151488178294e-14 K=2.62 tau=9.304724675465606e-08 off=-0.1

*Grain_516:
XU_516 in out fe_tanh Vc=0.2580964020134296 Qo=1.5673642828977376e-13 K=2.62 tau=1.0538488918950261e-07 off=-0.1

*Grain_517:
XU_517 in out fe_tanh Vc=0.7946175003565761 Qo=6.761747882026619e-13 K=2.62 tau=8.638966567418543e-08 off=-0.1

*Grain_518:
XU_518 in out fe_tanh Vc=0.10596299976245993 Qo=4.926675162301058e-14 K=2.62 tau=1.1473267285974081e-07 off=-0.1

*Grain_519:
XU_519 in out fe_tanh Vc=0.711127617095539 Qo=5.853090228211027e-13 K=2.62 tau=9.789591408996664e-08 off=-0.1

*Grain_520:
XU_520 in out fe_tanh Vc=0.42262539412671096 Qo=2.975744748555567e-13 K=2.62 tau=9.337551864616077e-08 off=-0.1

*Grain_521:
XU_521 in out fe_tanh Vc=0.8874380212952024 Qo=7.8060773715852e-13 K=2.62 tau=1.0426942448098339e-07 off=-0.1

*Grain_522:
XU_522 in out fe_tanh Vc=0.3069293991711135 Qo=1.9633758575617111e-13 K=2.62 tau=8.602353032946259e-08 off=-0.1

*Grain_523:
XU_523 in out fe_tanh Vc=0.4165420548094211 Qo=2.9201820160939406e-13 K=2.62 tau=9.98621475760137e-08 off=-0.1

*Grain_524:
XU_524 in out fe_tanh Vc=0.52289657815601 Qo=3.9245869028004925e-13 K=2.62 tau=9.303236407992647e-08 off=-0.1

*Grain_525:
XU_525 in out fe_tanh Vc=0.20159812735638838 Qo=1.1368046782413837e-13 K=2.62 tau=9.392157694791429e-08 off=-0.1

*Grain_526:
XU_526 in out fe_tanh Vc=0.3660838204543651 Qo=2.468926186744555e-13 K=2.62 tau=1.0429943343419398e-07 off=-0.1

*Grain_527:
XU_527 in out fe_tanh Vc=0.5231489666294009 Qo=3.9270496648813285e-13 K=2.62 tau=1.0261893443151421e-07 off=-0.1

*Grain_528:
XU_528 in out fe_tanh Vc=-0.05011288100521316 Qo=1.8611766399780337e-14 K=2.62 tau=8.591745322822849e-08 off=-0.1

*Grain_529:
XU_529 in out fe_tanh Vc=0.23940405683125968 Qo=1.4214263681858349e-13 K=2.62 tau=1.1793030397359822e-07 off=-0.1

*Grain_530:
XU_530 in out fe_tanh Vc=0.4634092245379728 Qo=3.354343137305329e-13 K=2.62 tau=9.044269786734624e-08 off=-0.1

*Grain_531:
XU_531 in out fe_tanh Vc=0.7606314985268579 Qo=6.38822212020767e-13 K=2.62 tau=9.435100212472628e-08 off=-0.1

*Grain_532:
XU_532 in out fe_tanh Vc=-0.08476897230048702 Qo=3.6860515435311474e-14 K=2.62 tau=1.1299149581941994e-07 off=-0.1

*Grain_533:
XU_533 in out fe_tanh Vc=0.09662131232295962 Qo=4.3696657920297087e-14 K=2.62 tau=1.2867095261211443e-07 off=-0.1

*Grain_534:
XU_534 in out fe_tanh Vc=-0.09796841140575863 Qo=4.4490296089226024e-14 K=2.62 tau=7.279277455837632e-08 off=-0.1

*Grain_535:
XU_535 in out fe_tanh Vc=0.8333772711058447 Qo=7.193621075615066e-13 K=2.62 tau=6.825914290722854e-08 off=-0.1

*Grain_536:
XU_536 in out fe_tanh Vc=0.48479428905577626 Qo=3.556953224930581e-13 K=2.62 tau=9.127532232774699e-08 off=-0.1

*Grain_537:
XU_537 in out fe_tanh Vc=0.4219162181225455 Qo=2.969254996547115e-13 K=2.62 tau=1.107244889769579e-07 off=-0.1

*Grain_538:
XU_538 in out fe_tanh Vc=0.701811883289958 Qo=5.753608975963692e-13 K=2.62 tau=9.744451459646839e-08 off=-0.1

*Grain_539:
XU_539 in out fe_tanh Vc=0.558393086872297 Qo=4.274402874315366e-13 K=2.62 tau=1.1574022517218372e-07 off=-0.1

*Grain_540:
XU_540 in out fe_tanh Vc=0.96356934697909 Qo=8.687629252165382e-13 K=2.62 tau=1.2403790848781665e-07 off=-0.1

*Grain_541:
XU_541 in out fe_tanh Vc=0.38621469061216307 Qo=2.6468591806543855e-13 K=2.62 tau=7.410861207470468e-08 off=-0.1

*Grain_542:
XU_542 in out fe_tanh Vc=0.5046861691771684 Qo=3.7478416610896586e-13 K=2.62 tau=1.0471388262012765e-07 off=-0.1

*Grain_543:
XU_543 in out fe_tanh Vc=0.4727256445653939 Qo=3.4422730912076884e-13 K=2.62 tau=9.351222959964891e-08 off=-0.1

*Grain_544:
XU_544 in out fe_tanh Vc=0.778457297844936 Qo=6.583527335678501e-13 K=2.62 tau=1.207547525393197e-07 off=-0.1

*Grain_545:
XU_545 in out fe_tanh Vc=0.6497870944330599 Qo=5.205420479209392e-13 K=2.62 tau=1.0159813426958672e-07 off=-0.1

*Grain_546:
XU_546 in out fe_tanh Vc=0.537480500004889 Qo=4.067475415697114e-13 K=2.62 tau=1.1890822920905611e-07 off=-0.1

*Grain_547:
XU_547 in out fe_tanh Vc=0.7796550576497099 Qo=6.596698892845684e-13 K=2.62 tau=1.0011669709604781e-07 off=-0.1

*Grain_548:
XU_548 in out fe_tanh Vc=0.33910038778072654 Qo=2.2350136649968962e-13 K=2.62 tau=9.492672175793904e-08 off=-0.1

*Grain_549:
XU_549 in out fe_tanh Vc=0.7123225901384413 Qo=5.865879580358354e-13 K=2.62 tau=9.393721510620547e-08 off=-0.1

*Grain_550:
XU_550 in out fe_tanh Vc=0.3510445507556401 Qo=2.3378913122422105e-13 K=2.62 tau=1.0381543866717575e-07 off=-0.1

*Grain_551:
XU_551 in out fe_tanh Vc=0.32906050768718653 Qo=2.1493735633068975e-13 K=2.62 tau=1.1038125710388218e-07 off=-0.1

*Grain_552:
XU_552 in out fe_tanh Vc=0.5329201242177632 Qo=4.0226677803400783e-13 K=2.62 tau=1.0158211991504012e-07 off=-0.1

*Grain_553:
XU_553 in out fe_tanh Vc=0.489566110644995 Qo=3.6025346065182076e-13 K=2.62 tau=1.1113362750798933e-07 off=-0.1

*Grain_554:
XU_554 in out fe_tanh Vc=0.23694416313092925 Qo=1.4024688682594169e-13 K=2.62 tau=9.784482551494071e-08 off=-0.1

*Grain_555:
XU_555 in out fe_tanh Vc=0.23086810082056952 Qo=1.3558964381629297e-13 K=2.62 tau=9.199038938474862e-08 off=-0.1

*Grain_556:
XU_556 in out fe_tanh Vc=0.12641039219852868 Qo=6.196850556677817e-14 K=2.62 tau=8.587021019084704e-08 off=-0.1

*Grain_557:
XU_557 in out fe_tanh Vc=0.5365414230576171 Qo=4.058239225325133e-13 K=2.62 tau=9.92283342068398e-08 off=-0.1

*Grain_558:
XU_558 in out fe_tanh Vc=0.837577652324486 Qo=7.240791066921864e-13 K=2.62 tau=1.020794615381781e-07 off=-0.1

*Grain_559:
XU_559 in out fe_tanh Vc=0.6744535007813361 Qo=5.463752618580316e-13 K=2.62 tau=1.1055101792776035e-07 off=-0.1

*Grain_560:
XU_560 in out fe_tanh Vc=0.548085169493117 Qo=4.1721112113811863e-13 K=2.62 tau=1.1194450217788462e-07 off=-0.1

*Grain_561:
XU_561 in out fe_tanh Vc=0.8131133368819201 Qo=6.967064325651555e-13 K=2.62 tau=1.1792250725211025e-07 off=-0.1

*Grain_562:
XU_562 in out fe_tanh Vc=0.4134868338122458 Qo=2.8923683555090366e-13 K=2.62 tau=1.1058359520074126e-07 off=-0.1

*Grain_563:
XU_563 in out fe_tanh Vc=0.23389407842612828 Qo=1.3790448959856488e-13 K=2.62 tau=1.0287215874690287e-07 off=-0.1

*Grain_564:
XU_564 in out fe_tanh Vc=1.097177683204122 Qo=1.0285217153100892e-12 K=2.62 tau=9.452562680223663e-08 off=-0.1

*Grain_565:
XU_565 in out fe_tanh Vc=0.15875084893051838 Qo=8.332671937872701e-14 K=2.62 tau=1.077523348934998e-07 off=-0.1

*Grain_566:
XU_566 in out fe_tanh Vc=0.6131416072532304 Qo=4.827057084537138e-13 K=2.62 tau=1.055814390800058e-07 off=-0.1

*Grain_567:
XU_567 in out fe_tanh Vc=0.44123333141019955 Qo=3.1471845919486705e-13 K=2.62 tau=9.664002546507278e-08 off=-0.1

*Grain_568:
XU_568 in out fe_tanh Vc=0.5197301624474314 Qo=3.893719917649699e-13 K=2.62 tau=9.661619476410363e-08 off=-0.1

*Grain_569:
XU_569 in out fe_tanh Vc=0.9675280061245939 Qo=8.734056940437839e-13 K=2.62 tau=8.793596546176907e-08 off=-0.1

*Grain_570:
XU_570 in out fe_tanh Vc=0.7988864482454172 Qo=6.809010138383377e-13 K=2.62 tau=1.0876148406103216e-07 off=-0.1

*Grain_571:
XU_571 in out fe_tanh Vc=0.3343994146564271 Qo=2.19481829473042e-13 K=2.62 tau=9.46965658156621e-08 off=-0.1

*Grain_572:
XU_572 in out fe_tanh Vc=0.7430051853259345 Qo=6.196447985541201e-13 K=2.62 tau=9.142312818443187e-08 off=-0.1

*Grain_573:
XU_573 in out fe_tanh Vc=0.6660181455039578 Qo=5.375084431169261e-13 K=2.62 tau=1.0879353239195105e-07 off=-0.1

*Grain_574:
XU_574 in out fe_tanh Vc=0.6902120896237622 Qo=5.630289694074077e-13 K=2.62 tau=1.0004903987604361e-07 off=-0.1

*Grain_575:
XU_575 in out fe_tanh Vc=0.058306622091321036 Qo=2.2661395840587764e-14 K=2.62 tau=1.0999248589429329e-07 off=-0.1

*Grain_576:
XU_576 in out fe_tanh Vc=0.7107234413338737 Qo=5.848765943701889e-13 K=2.62 tau=1.1349227869290672e-07 off=-0.1

*Grain_577:
XU_577 in out fe_tanh Vc=1.0405385415402777 Qo=9.600393470165706e-13 K=2.62 tau=9.952580799665797e-08 off=-0.1

*Grain_578:
XU_578 in out fe_tanh Vc=-0.07182931203105125 Qo=2.9719782675514966e-14 K=2.62 tau=8.921806402532661e-08 off=-0.1

*Grain_579:
XU_579 in out fe_tanh Vc=0.3265031487845833 Qo=2.127683357388085e-13 K=2.62 tau=8.73578055396527e-08 off=-0.1

*Grain_580:
XU_580 in out fe_tanh Vc=-0.06235024837622716 Qo=2.4725384539298132e-14 K=2.62 tau=9.968493150310394e-08 off=-0.1

*Grain_581:
XU_581 in out fe_tanh Vc=0.4442926028784668 Qo=3.175581168442212e-13 K=2.62 tau=1.0966192168889708e-07 off=-0.1

*Grain_582:
XU_582 in out fe_tanh Vc=0.5097708461346353 Qo=3.797002676368018e-13 K=2.62 tau=9.589777883999893e-08 off=-0.1

*Grain_583:
XU_583 in out fe_tanh Vc=0.6668720003219593 Qo=5.38404447426028e-13 K=2.62 tau=1.2162610544404145e-07 off=-0.1

*Grain_584:
XU_584 in out fe_tanh Vc=0.3408640854811774 Qo=2.2501373518754738e-13 K=2.62 tau=1.0939196758510779e-07 off=-0.1

*Grain_585:
XU_585 in out fe_tanh Vc=0.4400602123651698 Qo=3.1363111760662736e-13 K=2.62 tau=7.037057618541616e-08 off=-0.1

*Grain_586:
XU_586 in out fe_tanh Vc=0.8594414779135031 Qo=7.487461681890231e-13 K=2.62 tau=8.275197949319673e-08 off=-0.1

*Grain_587:
XU_587 in out fe_tanh Vc=0.8924502937583205 Qo=7.863441465736851e-13 K=2.62 tau=9.702389357628882e-08 off=-0.1

*Grain_588:
XU_588 in out fe_tanh Vc=0.6895386309224939 Qo=5.623149024817542e-13 K=2.62 tau=1.0362358207290184e-07 off=-0.1

*Grain_589:
XU_589 in out fe_tanh Vc=0.7102370030410917 Qo=5.843562508934604e-13 K=2.62 tau=9.896220908371609e-08 off=-0.1

*Grain_590:
XU_590 in out fe_tanh Vc=0.4313564301644583 Qo=3.055910071079018e-13 K=2.62 tau=9.650939472304035e-08 off=-0.1

*Grain_591:
XU_591 in out fe_tanh Vc=-0.20029526485232085 Qo=1.1272631168391525e-13 K=2.62 tau=8.425722461292482e-08 off=-0.1

*Grain_592:
XU_592 in out fe_tanh Vc=0.18696125521690313 Qo=1.0306958090036229e-13 K=2.62 tau=9.138184914231694e-08 off=-0.1

*Grain_593:
XU_593 in out fe_tanh Vc=0.6824568131327885 Qo=5.548187586960253e-13 K=2.62 tau=9.926198809007408e-08 off=-0.1

*Grain_594:
XU_594 in out fe_tanh Vc=0.4574436008481104 Qo=3.298315791598827e-13 K=2.62 tau=1.1393244404084377e-07 off=-0.1

*Grain_595:
XU_595 in out fe_tanh Vc=0.5067282579589488 Qo=3.767567753571006e-13 K=2.62 tau=9.591664009988929e-08 off=-0.1

*Grain_596:
XU_596 in out fe_tanh Vc=0.4727109881583285 Qo=3.4421343501470225e-13 K=2.62 tau=1.0699927936632138e-07 off=-0.1

*Grain_597:
XU_597 in out fe_tanh Vc=1.0630634977398712 Qo=9.871437004187334e-13 K=2.62 tau=1.1161345582217083e-07 off=-0.1

*Grain_598:
XU_598 in out fe_tanh Vc=0.4971459642453095 Qo=3.6752129160956563e-13 K=2.62 tau=8.810502787734099e-08 off=-0.1

*Grain_599:
XU_599 in out fe_tanh Vc=0.4305719169819491 Qo=3.0486868759644196e-13 K=2.62 tau=1.0800630585983544e-07 off=-0.1

*Grain_600:
XU_600 in out fe_tanh Vc=0.5112057644677795 Qo=3.8109028317906133e-13 K=2.62 tau=1.1458564152791424e-07 off=-0.1

*Grain_601:
XU_601 in out fe_tanh Vc=0.5633706016789126 Qo=4.324001590883818e-13 K=2.62 tau=8.662358829016352e-08 off=-0.1

*Grain_602:
XU_602 in out fe_tanh Vc=0.42341513676685116 Qo=2.982975620805599e-13 K=2.62 tau=9.724928006124131e-08 off=-0.1

*Grain_603:
XU_603 in out fe_tanh Vc=0.2773638379794652 Qo=1.7211479347027651e-13 K=2.62 tau=9.992475928780633e-08 off=-0.1

*Grain_604:
XU_604 in out fe_tanh Vc=0.11008786770173579 Qo=5.177435632815345e-14 K=2.62 tau=1.0340839479801726e-07 off=-0.1

*Grain_605:
XU_605 in out fe_tanh Vc=0.2628189610773831 Qo=1.6047489969147041e-13 K=2.62 tau=9.554985479285041e-08 off=-0.1

*Grain_606:
XU_606 in out fe_tanh Vc=0.2516037439544114 Qo=1.5163017614942752e-13 K=2.62 tau=1.0295864566189203e-07 off=-0.1

*Grain_607:
XU_607 in out fe_tanh Vc=0.20831929021846177 Qo=1.1863197038432678e-13 K=2.62 tau=1.0326944695122995e-07 off=-0.1

*Grain_608:
XU_608 in out fe_tanh Vc=0.22234851878152004 Qo=1.2912130992591896e-13 K=2.62 tau=1.0687777871637101e-07 off=-0.1

*Grain_609:
XU_609 in out fe_tanh Vc=-0.00955203411516925 Qo=2.157635280073648e-15 K=2.62 tau=9.691887121439327e-08 off=-0.1

*Grain_610:
XU_610 in out fe_tanh Vc=0.7723703650794725 Qo=6.516684464510671e-13 K=2.62 tau=1.0799831482016301e-07 off=-0.1

*Grain_611:
XU_611 in out fe_tanh Vc=0.17359988020898653 Qo=9.359823471960126e-14 K=2.62 tau=1.0967616606156662e-07 off=-0.1

*Grain_612:
XU_612 in out fe_tanh Vc=0.5913184821551365 Qo=4.604911625537557e-13 K=2.62 tau=1.2410942824416025e-07 off=-0.1

*Grain_613:
XU_613 in out fe_tanh Vc=0.41134994277823483 Qo=2.8729514309257894e-13 K=2.62 tau=1.1143875207503597e-07 off=-0.1

*Grain_614:
XU_614 in out fe_tanh Vc=0.31477466906509455 Qo=2.0288648554757251e-13 K=2.62 tau=1.0154657838748854e-07 off=-0.1

*Grain_615:
XU_615 in out fe_tanh Vc=0.2111090014439622 Qo=1.2070136663569067e-13 K=2.62 tau=1.0255653079035771e-07 off=-0.1

*Grain_616:
XU_616 in out fe_tanh Vc=0.46566849836331936 Qo=3.3756182641986655e-13 K=2.62 tau=1.0087778536915236e-07 off=-0.1

*Grain_617:
XU_617 in out fe_tanh Vc=0.7579083444930897 Qo=6.358506296018647e-13 K=2.62 tau=9.92324974110311e-08 off=-0.1

*Grain_618:
XU_618 in out fe_tanh Vc=0.40284720414142144 Qo=2.795991652480325e-13 K=2.62 tau=1.2477442998714434e-07 off=-0.1

*Grain_619:
XU_619 in out fe_tanh Vc=0.3663225038928031 Qo=2.471019025040868e-13 K=2.62 tau=1.1605842065432698e-07 off=-0.1

*Grain_620:
XU_620 in out fe_tanh Vc=0.5392832227328681 Qo=4.0852194668253846e-13 K=2.62 tau=1.0598948742283794e-07 off=-0.1

*Grain_621:
XU_621 in out fe_tanh Vc=1.0550767710744633 Qo=9.775133345997744e-13 K=2.62 tau=1.1518200159237573e-07 off=-0.1

*Grain_622:
XU_622 in out fe_tanh Vc=-0.1642134038801979 Qo=8.707321794353816e-14 K=2.62 tau=9.86095702498977e-08 off=-0.1

*Grain_623:
XU_623 in out fe_tanh Vc=0.23138723397240132 Qo=1.3598613276634931e-13 K=2.62 tau=1.0109005747456963e-07 off=-0.1

*Grain_624:
XU_624 in out fe_tanh Vc=0.4492152858686876 Qo=3.221397328689558e-13 K=2.62 tau=1.0240682078030359e-07 off=-0.1

*Grain_625:
XU_625 in out fe_tanh Vc=0.33700737742682113 Qo=2.217096727762477e-13 K=2.62 tau=1.1055427418815872e-07 off=-0.1

*Grain_626:
XU_626 in out fe_tanh Vc=-0.04651913973151123 Qo=1.6895637680206766e-14 K=2.62 tau=1.0422583270870389e-07 off=-0.1

*Grain_627:
XU_627 in out fe_tanh Vc=0.5338879725291636 Qo=4.032167722020099e-13 K=2.62 tau=1.1463185274578643e-07 off=-0.1

*Grain_628:
XU_628 in out fe_tanh Vc=-0.6970070287372231 Qo=5.702453011263382e-13 K=2.62 tau=9.618727594704305e-08 off=-0.1

*Grain_629:
XU_629 in out fe_tanh Vc=0.7009352808660995 Qo=5.74426817226899e-13 K=2.62 tau=9.22186386672445e-08 off=-0.1

*Grain_630:
XU_630 in out fe_tanh Vc=0.36190275496355173 Qo=2.4323320721198005e-13 K=2.62 tau=1.0296858918743888e-07 off=-0.1

*Grain_631:
XU_631 in out fe_tanh Vc=0.7309957358839254 Qo=6.066562931421585e-13 K=2.62 tau=9.685107312535788e-08 off=-0.1

*Grain_632:
XU_632 in out fe_tanh Vc=0.48460704563258955 Qo=3.555167373114456e-13 K=2.62 tau=1.0978055418216067e-07 off=-0.1

*Grain_633:
XU_633 in out fe_tanh Vc=0.8205795404646912 Qo=7.050343881250773e-13 K=2.62 tau=1.0800665958347869e-07 off=-0.1

*Grain_634:
XU_634 in out fe_tanh Vc=-0.35730161874055166 Qo=2.3922077295904953e-13 K=2.62 tau=1.1951201198859937e-07 off=-0.1

*Grain_635:
XU_635 in out fe_tanh Vc=0.129817027150537 Qo=6.414821375536992e-14 K=2.62 tau=9.769134678115956e-08 off=-0.1

*Grain_636:
XU_636 in out fe_tanh Vc=0.3876239816657935 Qo=2.6594218965246807e-13 K=2.62 tau=8.27105546262544e-08 off=-0.1

*Grain_637:
XU_637 in out fe_tanh Vc=0.10168694403725043 Qo=4.6697987545830476e-14 K=2.62 tau=1.1215932071200512e-07 off=-0.1

*Grain_638:
XU_638 in out fe_tanh Vc=0.5884805350693112 Qo=4.576201547115309e-13 K=2.62 tau=1.0691325489923695e-07 off=-0.1

*Grain_639:
XU_639 in out fe_tanh Vc=-0.05903631977546969 Qo=2.303077061738318e-14 K=2.62 tau=1.0502590726287188e-07 off=-0.1

*Grain_640:
XU_640 in out fe_tanh Vc=0.39011947482737735 Qo=2.68170085589166e-13 K=2.62 tau=9.98531225957828e-08 off=-0.1

*Grain_641:
XU_641 in out fe_tanh Vc=-0.010815235180861915 Qo=2.5357134165434116e-15 K=2.62 tau=9.460882272710806e-08 off=-0.1

*Grain_642:
XU_642 in out fe_tanh Vc=-0.37435061763710376 Qo=2.541648742782858e-13 K=2.62 tau=9.142082552815486e-08 off=-0.1

*Grain_643:
XU_643 in out fe_tanh Vc=0.5025597775512619 Qo=3.7273266569897606e-13 K=2.62 tau=1.0072551526020094e-07 off=-0.1

*Grain_644:
XU_644 in out fe_tanh Vc=-0.22201466832553562 Qo=1.2886933278079994e-13 K=2.62 tau=1.0747794709851225e-07 off=-0.1

*Grain_645:
XU_645 in out fe_tanh Vc=0.8207012982269972 Qo=7.051703882451109e-13 K=2.62 tau=1.0174741655561338e-07 off=-0.1

*Grain_646:
XU_646 in out fe_tanh Vc=0.27111471053738345 Qo=1.670907537264446e-13 K=2.62 tau=9.117981622190727e-08 off=-0.1

*Grain_647:
XU_647 in out fe_tanh Vc=0.6100312220313662 Qo=4.795248218054142e-13 K=2.62 tau=8.958420726378832e-08 off=-0.1

*Grain_648:
XU_648 in out fe_tanh Vc=0.2781649330051514 Qo=1.7276131610527855e-13 K=2.62 tau=1.0380950364122681e-07 off=-0.1

*Grain_649:
XU_649 in out fe_tanh Vc=0.5577262277452628 Qo=4.2677679641764363e-13 K=2.62 tau=8.42439063618297e-08 off=-0.1

*Grain_650:
XU_650 in out fe_tanh Vc=0.09776275611336666 Qo=4.4368922097968733e-14 K=2.62 tau=1.2252348800303456e-07 off=-0.1

*Grain_651:
XU_651 in out fe_tanh Vc=-0.029254531583918608 Qo=9.244948659913775e-15 K=2.62 tau=9.239722306685508e-08 off=-0.1

*Grain_652:
XU_652 in out fe_tanh Vc=0.6369418355707568 Qo=5.072045234404355e-13 K=2.62 tau=1.0165161042500825e-07 off=-0.1

*Grain_653:
XU_653 in out fe_tanh Vc=-0.30115921432382975 Qo=1.9155275938832307e-13 K=2.62 tau=1.1360242142983493e-07 off=-0.1

*Grain_654:
XU_654 in out fe_tanh Vc=-0.1626204729070576 Qo=8.597678398132445e-14 K=2.62 tau=8.745810976625257e-08 off=-0.1

*Grain_655:
XU_655 in out fe_tanh Vc=0.3171208253670533 Qo=2.048545443655992e-13 K=2.62 tau=1.0323519914899176e-07 off=-0.1

*Grain_656:
XU_656 in out fe_tanh Vc=0.32040712359508433 Qo=2.076185829511702e-13 K=2.62 tau=1.1383247544368701e-07 off=-0.1

*Grain_657:
XU_657 in out fe_tanh Vc=0.4940039722999479 Qo=3.6450457519828896e-13 K=2.62 tau=1.1716525160948052e-07 off=-0.1

*Grain_658:
XU_658 in out fe_tanh Vc=0.45862932147302193 Qo=3.3094343665155535e-13 K=2.62 tau=1.0284223566870982e-07 off=-0.1

*Grain_659:
XU_659 in out fe_tanh Vc=-0.26277046495798373 Qo=1.604364060729548e-13 K=2.62 tau=8.717928200633485e-08 off=-0.1

*Grain_660:
XU_660 in out fe_tanh Vc=0.3994658514381457 Qo=2.7655210440995533e-13 K=2.62 tau=9.713831814998191e-08 off=-0.1

*Grain_661:
XU_661 in out fe_tanh Vc=0.13848705753798535 Qo=6.97726719439793e-14 K=2.62 tau=1.1023226620289147e-07 off=-0.1

*Grain_662:
XU_662 in out fe_tanh Vc=0.19666545526668958 Qo=1.1007784449655958e-13 K=2.62 tau=1.0282444665568197e-07 off=-0.1

*Grain_663:
XU_663 in out fe_tanh Vc=0.35691169652479404 Qo=2.3888144931521034e-13 K=2.62 tau=8.787023240337186e-08 off=-0.1

*Grain_664:
XU_664 in out fe_tanh Vc=0.2469107766963069 Qo=1.4796379775461243e-13 K=2.62 tau=9.835576692778945e-08 off=-0.1

*Grain_665:
XU_665 in out fe_tanh Vc=0.6367858555567744 Qo=5.070430579574835e-13 K=2.62 tau=9.661272679488765e-08 off=-0.1

*Grain_666:
XU_666 in out fe_tanh Vc=0.3849210576913716 Qo=2.635339563885468e-13 K=2.62 tau=7.427284593880791e-08 off=-0.1

*Grain_667:
XU_667 in out fe_tanh Vc=0.3324050465343005 Qo=2.1778165887701754e-13 K=2.62 tau=8.863260244707032e-08 off=-0.1

*Grain_668:
XU_668 in out fe_tanh Vc=0.9072945886615891 Qo=8.033896404027397e-13 K=2.62 tau=9.22365368946165e-08 off=-0.1

*Grain_669:
XU_669 in out fe_tanh Vc=0.39763218174295734 Qo=2.749029462333127e-13 K=2.62 tau=1.0071108036999739e-07 off=-0.1

*Grain_670:
XU_670 in out fe_tanh Vc=0.5667410299590341 Qo=4.3576612041997795e-13 K=2.62 tau=9.225483524245881e-08 off=-0.1

*Grain_671:
XU_671 in out fe_tanh Vc=-0.1806129308564901 Qo=9.854325480195477e-14 K=2.62 tau=1.0672199445045096e-07 off=-0.1

*Grain_672:
XU_672 in out fe_tanh Vc=0.1834641682706496 Qo=1.0057036902885418e-13 K=2.62 tau=9.617430956335473e-08 off=-0.1

*Grain_673:
XU_673 in out fe_tanh Vc=0.1851072895537916 Qo=1.0174287103134944e-13 K=2.62 tau=9.358913835951858e-08 off=-0.1

*Grain_674:
XU_674 in out fe_tanh Vc=0.7049481875248312 Qo=5.787057109070987e-13 K=2.62 tau=9.550532538332609e-08 off=-0.1

*Grain_675:
XU_675 in out fe_tanh Vc=0.7491911046747781 Qo=6.263596984549443e-13 K=2.62 tau=9.697220665361686e-08 off=-0.1

*Grain_676:
XU_676 in out fe_tanh Vc=0.05437153458842675 Qo=2.0693620409722123e-14 K=2.62 tau=1.2004795187834632e-07 off=-0.1

*Grain_677:
XU_677 in out fe_tanh Vc=0.698324131376053 Qo=5.716465347765512e-13 K=2.62 tau=1.0474106409501106e-07 off=-0.1

*Grain_678:
XU_678 in out fe_tanh Vc=-0.2251269945435277 Qo=1.3122278659636472e-13 K=2.62 tau=1.173207764975125e-07 off=-0.1

*Grain_679:
XU_679 in out fe_tanh Vc=0.5004772294182834 Qo=3.7072598703373997e-13 K=2.62 tau=1.0886576802962571e-07 off=-0.1

*Grain_680:
XU_680 in out fe_tanh Vc=0.11262635796662085 Qo=5.333170436196451e-14 K=2.62 tau=1.071586685652983e-07 off=-0.1

*Grain_681:
XU_681 in out fe_tanh Vc=0.14158513264260436 Qo=7.180858319404865e-14 K=2.62 tau=8.80571786012392e-08 off=-0.1

*Grain_682:
XU_682 in out fe_tanh Vc=0.44635966740477817 Qo=3.194801203252035e-13 K=2.62 tau=9.77673217491611e-08 off=-0.1

*Grain_683:
XU_683 in out fe_tanh Vc=0.07558678528794299 Qo=3.175653048633629e-14 K=2.62 tau=9.945765025803766e-08 off=-0.1

*Grain_684:
XU_684 in out fe_tanh Vc=0.46233986749414485 Qo=3.344284052567776e-13 K=2.62 tau=9.732172048281167e-08 off=-0.1

*Grain_685:
XU_685 in out fe_tanh Vc=0.6188343737757585 Qo=4.885400450931225e-13 K=2.62 tau=1.0651527413194767e-07 off=-0.1

*Grain_686:
XU_686 in out fe_tanh Vc=0.6737381707755212 Qo=5.456220455846786e-13 K=2.62 tau=9.792423259886935e-08 off=-0.1

*Grain_687:
XU_687 in out fe_tanh Vc=0.27528864331309966 Qo=1.704426173023575e-13 K=2.62 tau=1.172599154024472e-07 off=-0.1

*Grain_688:
XU_688 in out fe_tanh Vc=0.9668070928940892 Qo=8.725597721378521e-13 K=2.62 tau=9.593228739897977e-08 off=-0.1

*Grain_689:
XU_689 in out fe_tanh Vc=0.9261942278847446 Qo=8.252130770625874e-13 K=2.62 tau=1.0407631462511779e-07 off=-0.1

*Grain_690:
XU_690 in out fe_tanh Vc=0.373283262161313 Qo=2.5322319392935307e-13 K=2.62 tau=1.0121365915039682e-07 off=-0.1

*Grain_691:
XU_691 in out fe_tanh Vc=0.26847624702275685 Qo=1.6497990120024395e-13 K=2.62 tau=1.1126273163250376e-07 off=-0.1

*Grain_692:
XU_692 in out fe_tanh Vc=0.31365648620274444 Qo=2.019500500676066e-13 K=2.62 tau=9.260705438039073e-08 off=-0.1

*Grain_693:
XU_693 in out fe_tanh Vc=0.26766003323311877 Qo=1.6432816144134558e-13 K=2.62 tau=1.0444036267162313e-07 off=-0.1

*Grain_694:
XU_694 in out fe_tanh Vc=0.4174372551394472 Qo=2.928343226282701e-13 K=2.62 tau=1.0012823340896958e-07 off=-0.1

*Grain_695:
XU_695 in out fe_tanh Vc=0.32875069297393417 Qo=2.146743173101913e-13 K=2.62 tau=1.0503032338379896e-07 off=-0.1

*Grain_696:
XU_696 in out fe_tanh Vc=0.4262474449796127 Qo=3.008941441551898e-13 K=2.62 tau=1.0583424537621434e-07 off=-0.1

*Grain_697:
XU_697 in out fe_tanh Vc=0.2938862985618569 Qo=1.8556093459063868e-13 K=2.62 tau=9.219445387783324e-08 off=-0.1

*Grain_698:
XU_698 in out fe_tanh Vc=0.09361420083043426 Qo=4.193702947325652e-14 K=2.62 tau=9.699178071737889e-08 off=-0.1

*Grain_699:
XU_699 in out fe_tanh Vc=0.4164807258347634 Qo=2.9196230949602123e-13 K=2.62 tau=1.1919299354069972e-07 off=-0.1

*Grain_700:
XU_700 in out fe_tanh Vc=0.38046232849293593 Qo=2.595724345563335e-13 K=2.62 tau=1.0395251379136963e-07 off=-0.1

*Grain_701:
XU_701 in out fe_tanh Vc=-0.17276528010469572 Qo=9.301367838542456e-14 K=2.62 tau=9.089285457214678e-08 off=-0.1

*Grain_702:
XU_702 in out fe_tanh Vc=0.9184076948350307 Qo=8.162056154164224e-13 K=2.62 tau=1.105700159203534e-07 off=-0.1

*Grain_703:
XU_703 in out fe_tanh Vc=0.599049547776796 Qo=4.683332351575061e-13 K=2.62 tau=8.808656842874119e-08 off=-0.1

*Grain_704:
XU_704 in out fe_tanh Vc=0.27401893373708164 Qo=1.694213562850181e-13 K=2.62 tau=1.0738774252932391e-07 off=-0.1

*Grain_705:
XU_705 in out fe_tanh Vc=0.33043805632679224 Qo=2.1610782231316162e-13 K=2.62 tau=1.1005508940061226e-07 off=-0.1

*Grain_706:
XU_706 in out fe_tanh Vc=0.2673103988292343 Qo=1.6404916359442545e-13 K=2.62 tau=1.1310136800567519e-07 off=-0.1

*Grain_707:
XU_707 in out fe_tanh Vc=0.8485152119122462 Qo=7.363951725797291e-13 K=2.62 tau=8.421661768231572e-08 off=-0.1

*Grain_708:
XU_708 in out fe_tanh Vc=0.42596829367568323 Qo=3.006379953771877e-13 K=2.62 tau=9.141760206941836e-08 off=-0.1

*Grain_709:
XU_709 in out fe_tanh Vc=0.38386227029966424 Qo=2.6259198506197524e-13 K=2.62 tau=9.045145028787628e-08 off=-0.1

*Grain_710:
XU_710 in out fe_tanh Vc=0.4966247474595894 Qo=3.6702045967680137e-13 K=2.62 tau=8.523011190537161e-08 off=-0.1

*Grain_711:
XU_711 in out fe_tanh Vc=0.5813025290210497 Qo=4.5037708591152664e-13 K=2.62 tau=9.074435803138316e-08 off=-0.1

*Grain_712:
XU_712 in out fe_tanh Vc=0.8093300045605174 Qo=6.924951630758871e-13 K=2.62 tau=7.134522425353168e-08 off=-0.1

*Grain_713:
XU_713 in out fe_tanh Vc=0.37950105801688017 Qo=2.587201764429275e-13 K=2.62 tau=1.1849450957035417e-07 off=-0.1

*Grain_714:
XU_714 in out fe_tanh Vc=0.9380120457830153 Qo=8.389273451979686e-13 K=2.62 tau=1.0139511809020295e-07 off=-0.1

*Grain_715:
XU_715 in out fe_tanh Vc=0.6947332873088197 Qo=5.678281919854346e-13 K=2.62 tau=1.2218937745385505e-07 off=-0.1

*Grain_716:
XU_716 in out fe_tanh Vc=0.3231329545492979 Qo=2.0991768945515175e-13 K=2.62 tau=8.188516108403739e-08 off=-0.1

*Grain_717:
XU_717 in out fe_tanh Vc=0.044773389798200613 Qo=1.6076051151340362e-14 K=2.62 tau=9.60607334940876e-08 off=-0.1

*Grain_718:
XU_718 in out fe_tanh Vc=0.40540699375849104 Qo=2.819109972722239e-13 K=2.62 tau=8.869621177516184e-08 off=-0.1

*Grain_719:
XU_719 in out fe_tanh Vc=0.03947728560365815 Qo=1.3649127138302758e-14 K=2.62 tau=1.0944296368572953e-07 off=-0.1

*Grain_720:
XU_720 in out fe_tanh Vc=0.11269919785004123 Qo=5.337654792786336e-14 K=2.62 tau=1.1058774003949036e-07 off=-0.1

*Grain_721:
XU_721 in out fe_tanh Vc=0.8530360533560364 Qo=7.414997576253226e-13 K=2.62 tau=8.931349463388795e-08 off=-0.1

*Grain_722:
XU_722 in out fe_tanh Vc=0.7278998027457457 Qo=6.033182916441179e-13 K=2.62 tau=9.58091966076459e-08 off=-0.1

*Grain_723:
XU_723 in out fe_tanh Vc=0.4792884057814914 Qo=3.504527003857693e-13 K=2.62 tau=8.911852447138839e-08 off=-0.1

*Grain_724:
XU_724 in out fe_tanh Vc=0.07857834080854531 Qo=3.3400050322004015e-14 K=2.62 tau=8.886798336964514e-08 off=-0.1

*Grain_725:
XU_725 in out fe_tanh Vc=0.4352434893042589 Qo=3.091757185311318e-13 K=2.62 tau=1.0629208467050956e-07 off=-0.1

*Grain_726:
XU_726 in out fe_tanh Vc=0.3829446691462176 Qo=2.617762530543828e-13 K=2.62 tau=1.0568512243402114e-07 off=-0.1

*Grain_727:
XU_727 in out fe_tanh Vc=0.4354301669909415 Qo=3.093481183459899e-13 K=2.62 tau=9.957464792458246e-08 off=-0.1

*Grain_728:
XU_728 in out fe_tanh Vc=0.7323341447917697 Qo=6.081006657448597e-13 K=2.62 tau=1.1351907039049937e-07 off=-0.1

*Grain_729:
XU_729 in out fe_tanh Vc=0.6361172926136143 Qo=5.063511175881464e-13 K=2.62 tau=9.541392815804869e-08 off=-0.1

*Grain_730:
XU_730 in out fe_tanh Vc=1.1647665966457144 Qo=1.1116395507357093e-12 K=2.62 tau=9.119592665477624e-08 off=-0.1

*Grain_731:
XU_731 in out fe_tanh Vc=0.14322574615499634 Qo=7.289216203499683e-14 K=2.62 tau=1.1087472155887357e-07 off=-0.1

*Grain_732:
XU_732 in out fe_tanh Vc=0.1384336016704295 Qo=6.973766213406439e-14 K=2.62 tau=1.0665317199670684e-07 off=-0.1

*Grain_733:
XU_733 in out fe_tanh Vc=0.23040199038877412 Qo=1.3523387886553182e-13 K=2.62 tau=1.0894996844699418e-07 off=-0.1

*Grain_734:
XU_734 in out fe_tanh Vc=0.07037270907347176 Qo=2.893869625538542e-14 K=2.62 tau=1.064105438598062e-07 off=-0.1

*Grain_735:
XU_735 in out fe_tanh Vc=0.49565852299388946 Qo=3.6609244150475803e-13 K=2.62 tau=9.636514632277583e-08 off=-0.1

*Grain_736:
XU_736 in out fe_tanh Vc=0.5398886774995011 Qo=4.0911829040302045e-13 K=2.62 tau=8.223886124408022e-08 off=-0.1

*Grain_737:
XU_737 in out fe_tanh Vc=0.05240443206696471 Qo=1.9725673242193722e-14 K=2.62 tau=1.0353260454452339e-07 off=-0.1

*Grain_738:
XU_738 in out fe_tanh Vc=0.4597327172258395 Qo=3.3197887257202065e-13 K=2.62 tau=1.0790506644006776e-07 off=-0.1

*Grain_739:
XU_739 in out fe_tanh Vc=0.4923872026066057 Qo=3.6295450760662716e-13 K=2.62 tau=9.363848792351997e-08 off=-0.1

*Grain_740:
XU_740 in out fe_tanh Vc=0.7461574528804003 Qo=6.230645410665589e-13 K=2.62 tau=1.1978693684673637e-07 off=-0.1

*Grain_741:
XU_741 in out fe_tanh Vc=0.43458217358895457 Qo=3.0856516146256784e-13 K=2.62 tau=1.1468146215936577e-07 off=-0.1

*Grain_742:
XU_742 in out fe_tanh Vc=0.5863361178720055 Qo=4.554535083941794e-13 K=2.62 tau=1.0086893711885333e-07 off=-0.1

*Grain_743:
XU_743 in out fe_tanh Vc=0.555794703273039 Qo=4.2485637098512344e-13 K=2.62 tau=9.05210267483166e-08 off=-0.1

*Grain_744:
XU_744 in out fe_tanh Vc=0.6750323617211096 Qo=5.469849566823662e-13 K=2.62 tau=1.0592664121117915e-07 off=-0.1

*Grain_745:
XU_745 in out fe_tanh Vc=0.5806891875429306 Qo=4.4975942373862435e-13 K=2.62 tau=9.338458913862556e-08 off=-0.1

*Grain_746:
XU_746 in out fe_tanh Vc=0.7972146379001921 Qo=6.790492189811577e-13 K=2.62 tau=8.209554271892213e-08 off=-0.1

*Grain_747:
XU_747 in out fe_tanh Vc=0.6041885889300465 Qo=4.735629144743576e-13 K=2.62 tau=1.0124252434860482e-07 off=-0.1

*Grain_748:
XU_748 in out fe_tanh Vc=0.9057845292050122 Qo=8.016518122532843e-13 K=2.62 tau=1.0430133670807832e-07 off=-0.1

*Grain_749:
XU_749 in out fe_tanh Vc=0.7942724450714242 Qo=6.757931036426113e-13 K=2.62 tau=1.0385957081011463e-07 off=-0.1

*Grain_750:
XU_750 in out fe_tanh Vc=0.8204263235830896 Qo=7.048632576236904e-13 K=2.62 tau=1.1261046151266969e-07 off=-0.1

*Grain_751:
XU_751 in out fe_tanh Vc=0.2857562891861326 Qo=1.7891549206886653e-13 K=2.62 tau=1.1738384083053903e-07 off=-0.1

*Grain_752:
XU_752 in out fe_tanh Vc=0.6600595857632248 Qo=5.312653552162001e-13 K=2.62 tau=1.1514995154523506e-07 off=-0.1

*Grain_753:
XU_753 in out fe_tanh Vc=0.3054522089471129 Qo=1.951100596360469e-13 K=2.62 tau=1.0188931926530967e-07 off=-0.1

*Grain_754:
XU_754 in out fe_tanh Vc=0.1638897503368568 Qo=8.685018385951785e-14 K=2.62 tau=9.466097990159162e-08 off=-0.1

*Grain_755:
XU_755 in out fe_tanh Vc=0.259466760643185 Qo=1.5781913518843505e-13 K=2.62 tau=1.010993748411759e-07 off=-0.1

*Grain_756:
XU_756 in out fe_tanh Vc=0.8383866502109892 Qo=7.249884221559662e-13 K=2.62 tau=7.429139176598956e-08 off=-0.1

*Grain_757:
XU_757 in out fe_tanh Vc=0.48276886453764567 Qo=3.5376465467830707e-13 K=2.62 tau=9.609604355491088e-08 off=-0.1

*Grain_758:
XU_758 in out fe_tanh Vc=0.5063013729465176 Qo=3.763442170718836e-13 K=2.62 tau=9.99198152573543e-08 off=-0.1

*Grain_759:
XU_759 in out fe_tanh Vc=0.13230601378400098 Qo=6.575168256713107e-14 K=2.62 tau=9.236213861710762e-08 off=-0.1

*Grain_760:
XU_760 in out fe_tanh Vc=0.6463584139540927 Qo=5.16974163311297e-13 K=2.62 tau=9.016842295008872e-08 off=-0.1

*Grain_761:
XU_761 in out fe_tanh Vc=0.3246716178547675 Qo=2.1121805207776839e-13 K=2.62 tau=9.0339973013032e-08 off=-0.1

*Grain_762:
XU_762 in out fe_tanh Vc=0.21008387929959038 Qo=1.1993997588686714e-13 K=2.62 tau=9.431826209388564e-08 off=-0.1

*Grain_763:
XU_763 in out fe_tanh Vc=-0.1833837427559173 Qo=1.0051305942221839e-13 K=2.62 tau=1.0660966950699516e-07 off=-0.1

*Grain_764:
XU_764 in out fe_tanh Vc=0.6930388593118946 Qo=5.660284663201352e-13 K=2.62 tau=8.800880086041119e-08 off=-0.1

*Grain_765:
XU_765 in out fe_tanh Vc=0.3988936929503512 Qo=2.7603727463324016e-13 K=2.62 tau=1.058219747043358e-07 off=-0.1

*Grain_766:
XU_766 in out fe_tanh Vc=0.6435289331855998 Qo=5.140340777305324e-13 K=2.62 tau=1.0293928741037256e-07 off=-0.1

*Grain_767:
XU_767 in out fe_tanh Vc=0.25027930333942644 Qo=1.505933620216775e-13 K=2.62 tau=1.0573074542399315e-07 off=-0.1

*Grain_768:
XU_768 in out fe_tanh Vc=0.01791799991399351 Qo=4.8879842701958554e-15 K=2.62 tau=9.716613949737288e-08 off=-0.1

*Grain_769:
XU_769 in out fe_tanh Vc=0.4203779222833019 Qo=2.9551891228776523e-13 K=2.62 tau=1.002996992361764e-07 off=-0.1

*Grain_770:
XU_770 in out fe_tanh Vc=0.6222154113784708 Qo=4.920128022355704e-13 K=2.62 tau=1.1029047318306846e-07 off=-0.1

*Grain_771:
XU_771 in out fe_tanh Vc=0.19179615747216772 Qo=1.0654799536209239e-13 K=2.62 tau=9.590512709800066e-08 off=-0.1

*Grain_772:
XU_772 in out fe_tanh Vc=1.102062233909968 Qo=1.0344782557445943e-12 K=2.62 tau=9.134076388431012e-08 off=-0.1

*Grain_773:
XU_773 in out fe_tanh Vc=0.10787484366924477 Qo=5.0425433862324916e-14 K=2.62 tau=1.0412501146202975e-07 off=-0.1

*Grain_774:
XU_774 in out fe_tanh Vc=0.4336407739292864 Qo=3.076964987871431e-13 K=2.62 tau=9.29247039734752e-08 off=-0.1

*Grain_775:
XU_775 in out fe_tanh Vc=0.819479915358265 Qo=7.038064109853618e-13 K=2.62 tau=1.2058306743013119e-07 off=-0.1

*Grain_776:
XU_776 in out fe_tanh Vc=0.4604123077663129 Qo=3.3261697730447694e-13 K=2.62 tau=1.2372958637228397e-07 off=-0.1

*Grain_777:
XU_777 in out fe_tanh Vc=0.5182964529216555 Qo=3.8797622950085957e-13 K=2.62 tau=9.24913823263733e-08 off=-0.1

*Grain_778:
XU_778 in out fe_tanh Vc=0.2957953279098549 Qo=1.871294380775853e-13 K=2.62 tau=1.0032231006324974e-07 off=-0.1

*Grain_779:
XU_779 in out fe_tanh Vc=0.06113030072115794 Qo=2.4098327507289205e-14 K=2.62 tau=1.0189652957310564e-07 off=-0.1

*Grain_780:
XU_780 in out fe_tanh Vc=0.8126186169115739 Qo=6.961554195120914e-13 K=2.62 tau=9.6349063925066e-08 off=-0.1

*Grain_781:
XU_781 in out fe_tanh Vc=0.7870287848191626 Qo=6.677919999244854e-13 K=2.62 tau=1.1216941750948199e-07 off=-0.1

*Grain_782:
XU_782 in out fe_tanh Vc=0.13555233035154995 Qo=6.785666246807286e-14 K=2.62 tau=9.99647946684234e-08 off=-0.1

*Grain_783:
XU_783 in out fe_tanh Vc=0.5322753487154459 Qo=4.0163418401634477e-13 K=2.62 tau=1.0602940674752789e-07 off=-0.1

*Grain_784:
XU_784 in out fe_tanh Vc=0.6157494107983167 Qo=4.853763560083681e-13 K=2.62 tau=9.074904593502436e-08 off=-0.1

*Grain_785:
XU_785 in out fe_tanh Vc=0.4796615328266062 Qo=3.5080741842186685e-13 K=2.62 tau=1.1641069623155148e-07 off=-0.1

*Grain_786:
XU_786 in out fe_tanh Vc=0.11268726873244955 Qo=5.336920322155837e-14 K=2.62 tau=1.0483858078432697e-07 off=-0.1

*Grain_787:
XU_787 in out fe_tanh Vc=0.5277132294771938 Qo=3.9716483294488213e-13 K=2.62 tau=9.213474287651925e-08 off=-0.1

*Grain_788:
XU_788 in out fe_tanh Vc=0.8089016248988126 Qo=6.920187004804332e-13 K=2.62 tau=9.302534799566403e-08 off=-0.1

*Grain_789:
XU_789 in out fe_tanh Vc=0.6272736220685471 Qo=4.972188022460687e-13 K=2.62 tau=1.0423377587046607e-07 off=-0.1

*Grain_790:
XU_790 in out fe_tanh Vc=0.45987046936580134 Qo=3.3210819273945606e-13 K=2.62 tau=8.078884974903416e-08 off=-0.1

*Grain_791:
XU_791 in out fe_tanh Vc=0.580586293338349 Qo=4.496558238579754e-13 K=2.62 tau=8.990502773300612e-08 off=-0.1

*Grain_792:
XU_792 in out fe_tanh Vc=0.12353599344177679 Qo=6.014298458730621e-14 K=2.62 tau=9.549615536964887e-08 off=-0.1

*Grain_793:
XU_793 in out fe_tanh Vc=0.46005783807165457 Qo=3.3228411103779123e-13 K=2.62 tau=9.04347906845408e-08 off=-0.1

*Grain_794:
XU_794 in out fe_tanh Vc=0.24908046582966437 Qo=1.49656291956547e-13 K=2.62 tau=9.304977084185394e-08 off=-0.1

*Grain_795:
XU_795 in out fe_tanh Vc=0.33852134263635086 Qo=2.2300534971303236e-13 K=2.62 tau=9.325224378072237e-08 off=-0.1

*Grain_796:
XU_796 in out fe_tanh Vc=0.5102958579953182 Qo=3.802087143525503e-13 K=2.62 tau=8.317938253195907e-08 off=-0.1

*Grain_797:
XU_797 in out fe_tanh Vc=0.33484765746342854 Qo=2.1986436962874928e-13 K=2.62 tau=1.0172313750643372e-07 off=-0.1

*Grain_798:
XU_798 in out fe_tanh Vc=0.8371418296642374 Qo=7.235893502108746e-13 K=2.62 tau=1.0430998390559825e-07 off=-0.1

*Grain_799:
XU_799 in out fe_tanh Vc=-0.015139967296428136 Qo=3.926592462729726e-15 K=2.62 tau=1.0931436806960518e-07 off=-0.1

*Grain_800:
XU_800 in out fe_tanh Vc=-0.262763487880022 Qo=1.6043086821803853e-13 K=2.62 tau=9.333146247427928e-08 off=-0.1

*Grain_801:
XU_801 in out fe_tanh Vc=0.6618305532393275 Qo=5.331191298323424e-13 K=2.62 tau=1.0917675181180847e-07 off=-0.1

*Grain_802:
XU_802 in out fe_tanh Vc=0.7111891972966269 Qo=5.853749140746749e-13 K=2.62 tau=9.720825069809251e-08 off=-0.1

*Grain_803:
XU_803 in out fe_tanh Vc=0.3962982396226424 Qo=2.7370466311727954e-13 K=2.62 tau=1.0350018439623794e-07 off=-0.1

*Grain_804:
XU_804 in out fe_tanh Vc=0.2889067880441812 Qo=1.8148405743261334e-13 K=2.62 tau=9.173632594683026e-08 off=-0.1

*Grain_805:
XU_805 in out fe_tanh Vc=-0.07402374790512511 Qo=3.0905501953356586e-14 K=2.62 tau=9.453162243624354e-08 off=-0.1

*Grain_806:
XU_806 in out fe_tanh Vc=0.3161262456090802 Qo=2.0401971195838288e-13 K=2.62 tau=1.0137822064795899e-07 off=-0.1

*Grain_807:
XU_807 in out fe_tanh Vc=0.6508834412867668 Qo=5.216841000256525e-13 K=2.62 tau=9.762813362045752e-08 off=-0.1

*Grain_808:
XU_808 in out fe_tanh Vc=0.4784676601715034 Qo=3.49672739552281e-13 K=2.62 tau=9.291583727885754e-08 off=-0.1

*Grain_809:
XU_809 in out fe_tanh Vc=0.1553262214406988 Qo=8.099750123385049e-14 K=2.62 tau=8.606657340739702e-08 off=-0.1

*Grain_810:
XU_810 in out fe_tanh Vc=0.978004973744764 Qo=8.857206965364547e-13 K=2.62 tau=7.950395042107374e-08 off=-0.1

*Grain_811:
XU_811 in out fe_tanh Vc=0.36828477082593364 Qo=2.488240181342715e-13 K=2.62 tau=9.948206133412348e-08 off=-0.1

*Grain_812:
XU_812 in out fe_tanh Vc=0.30790625192202525 Qo=1.9715031248337874e-13 K=2.62 tau=1.0489951877558906e-07 off=-0.1

*Grain_813:
XU_813 in out fe_tanh Vc=-0.1364363411603301 Qo=6.843251386321497e-14 K=2.62 tau=1.0037346436422599e-07 off=-0.1

*Grain_814:
XU_814 in out fe_tanh Vc=0.34920626494778617 Qo=2.3219883956695976e-13 K=2.62 tau=1.1295496948436384e-07 off=-0.1

*Grain_815:
XU_815 in out fe_tanh Vc=0.09530743948105252 Qo=4.292578569339831e-14 K=2.62 tau=1.0972857380813451e-07 off=-0.1

*Grain_816:
XU_816 in out fe_tanh Vc=0.34085926182556403 Qo=2.2500959570069076e-13 K=2.62 tau=9.2443340635899e-08 off=-0.1

*Grain_817:
XU_817 in out fe_tanh Vc=0.7710516657680417 Qo=6.502224109979463e-13 K=2.62 tau=1.0206431478821185e-07 off=-0.1

*Grain_818:
XU_818 in out fe_tanh Vc=0.3172042453460184 Qo=2.0492460134411864e-13 K=2.62 tau=1.0357725409519166e-07 off=-0.1

*Grain_819:
XU_819 in out fe_tanh Vc=1.1048188410281365 Qo=1.0378433427126342e-12 K=2.62 tau=1.0619237758839495e-07 off=-0.1

*Grain_820:
XU_820 in out fe_tanh Vc=0.597692330348046 Qo=4.669543207188546e-13 K=2.62 tau=1.0129138193702432e-07 off=-0.1

*Grain_821:
XU_821 in out fe_tanh Vc=0.6274696682178302 Qo=4.974208307020024e-13 K=2.62 tau=8.048064288619712e-08 off=-0.1

*Grain_822:
XU_822 in out fe_tanh Vc=0.3778851715904735 Qo=2.572889981217313e-13 K=2.62 tau=9.237232047119056e-08 off=-0.1

*Grain_823:
XU_823 in out fe_tanh Vc=0.24947149525459736 Qo=1.499617913291049e-13 K=2.62 tau=8.37989201951513e-08 off=-0.1

*Grain_824:
XU_824 in out fe_tanh Vc=0.896377847282107 Qo=7.908458863661505e-13 K=2.62 tau=1.089976401607721e-07 off=-0.1

*Grain_825:
XU_825 in out fe_tanh Vc=0.40004777170930567 Qo=2.770759448258496e-13 K=2.62 tau=1.1721732071109788e-07 off=-0.1

*Grain_826:
XU_826 in out fe_tanh Vc=0.6814142003527721 Qo=5.537171108515446e-13 K=2.62 tau=1.0018771687198695e-07 off=-0.1

*Grain_827:
XU_827 in out fe_tanh Vc=0.5094461141690453 Qo=3.793858602098739e-13 K=2.62 tau=1.1195062844004044e-07 off=-0.1

*Grain_828:
XU_828 in out fe_tanh Vc=0.2618258141204733 Qo=1.5968701832139144e-13 K=2.62 tau=7.97009505385428e-08 off=-0.1

*Grain_829:
XU_829 in out fe_tanh Vc=0.38848545256781997 Qo=2.667107982656437e-13 K=2.62 tau=7.567602832832067e-08 off=-0.1

*Grain_830:
XU_830 in out fe_tanh Vc=-0.06761359730643435 Qo=2.747246735233987e-14 K=2.62 tau=1.1608046485955954e-07 off=-0.1

*Grain_831:
XU_831 in out fe_tanh Vc=0.7683376824475079 Qo=6.472486953770396e-13 K=2.62 tau=1.0481913800981456e-07 off=-0.1

*Grain_832:
XU_832 in out fe_tanh Vc=0.6847570352743838 Qo=5.572510099457055e-13 K=2.62 tau=9.9782416088321e-08 off=-0.1

*Grain_833:
XU_833 in out fe_tanh Vc=0.48228374893845255 Qo=3.5330259475954976e-13 K=2.62 tau=8.621040596449899e-08 off=-0.1

*Grain_834:
XU_834 in out fe_tanh Vc=0.7231178912632523 Qo=5.981708557798294e-13 K=2.62 tau=9.699138920877486e-08 off=-0.1

*Grain_835:
XU_835 in out fe_tanh Vc=0.24825506652314586 Qo=1.4901190510766494e-13 K=2.62 tau=8.954134462613537e-08 off=-0.1

*Grain_836:
XU_836 in out fe_tanh Vc=0.6827029737249888 Qo=5.55078931164601e-13 K=2.62 tau=9.826558632335848e-08 off=-0.1

*Grain_837:
XU_837 in out fe_tanh Vc=0.6392672223901296 Qo=5.096130945174467e-13 K=2.62 tau=1.0000346075298045e-07 off=-0.1

*Grain_838:
XU_838 in out fe_tanh Vc=0.34859449507238904 Qo=2.3167015665724474e-13 K=2.62 tau=1.0919904105417014e-07 off=-0.1

*Grain_839:
XU_839 in out fe_tanh Vc=0.5960293776466381 Qo=4.652660637192969e-13 K=2.62 tau=1.0230554835642756e-07 off=-0.1

*Grain_840:
XU_840 in out fe_tanh Vc=0.5852285946450302 Qo=4.5433543457499984e-13 K=2.62 tau=1.0559738754056267e-07 off=-0.1

*Grain_841:
XU_841 in out fe_tanh Vc=0.5431436611307177 Qo=4.1232772746177813e-13 K=2.62 tau=8.665432854638705e-08 off=-0.1

*Grain_842:
XU_842 in out fe_tanh Vc=0.4859410903051813 Qo=3.5678954629559035e-13 K=2.62 tau=8.27933393740569e-08 off=-0.1

*Grain_843:
XU_843 in out fe_tanh Vc=0.7696611563171238 Qo=6.486984347240901e-13 K=2.62 tau=8.712356325304063e-08 off=-0.1

*Grain_844:
XU_844 in out fe_tanh Vc=0.08034019361284467 Qo=3.43768553425515e-14 K=2.62 tau=9.628286030735634e-08 off=-0.1

*Grain_845:
XU_845 in out fe_tanh Vc=0.3978680199804136 Qo=2.7511492583482536e-13 K=2.62 tau=1.0987282118243207e-07 off=-0.1

*Grain_846:
XU_846 in out fe_tanh Vc=0.4235421879557829 Qo=2.9841392777233513e-13 K=2.62 tau=8.051670630219888e-08 off=-0.1

*Grain_847:
XU_847 in out fe_tanh Vc=0.7008706748095327 Qo=5.743579888754583e-13 K=2.62 tau=1.020085155555545e-07 off=-0.1

*Grain_848:
XU_848 in out fe_tanh Vc=-0.11667099437980133 Qo=5.583482760903966e-14 K=2.62 tau=1.02933261493897e-07 off=-0.1

*Grain_849:
XU_849 in out fe_tanh Vc=0.2724804058032212 Qo=1.6818577898232504e-13 K=2.62 tau=9.47643140051295e-08 off=-0.1

*Grain_850:
XU_850 in out fe_tanh Vc=0.6102493772498587 Qo=4.797477634917212e-13 K=2.62 tau=9.756230575151817e-08 off=-0.1

*Grain_851:
XU_851 in out fe_tanh Vc=0.7126989229676 Qo=5.869908664105705e-13 K=2.62 tau=1.0630193157212716e-07 off=-0.1

*Grain_852:
XU_852 in out fe_tanh Vc=0.5863417214446496 Qo=4.554591669601818e-13 K=2.62 tau=1.1105335227693439e-07 off=-0.1

*Grain_853:
XU_853 in out fe_tanh Vc=0.39998362242728114 Qo=2.770181868888351e-13 K=2.62 tau=9.89882127734503e-08 off=-0.1

*Grain_854:
XU_854 in out fe_tanh Vc=0.3735509955871836 Qo=2.5345932744146167e-13 K=2.62 tau=1.1800873856114359e-07 off=-0.1

*Grain_855:
XU_855 in out fe_tanh Vc=0.5441119167334966 Qo=4.1328354999351994e-13 K=2.62 tau=1.0125485013041531e-07 off=-0.1

*Grain_856:
XU_856 in out fe_tanh Vc=0.03533294068204745 Qo=1.1816452948986623e-14 K=2.62 tau=1.0500121609278782e-07 off=-0.1

*Grain_857:
XU_857 in out fe_tanh Vc=0.3726013420471351 Qo=2.526219887062245e-13 K=2.62 tau=1.0453891828225806e-07 off=-0.1

*Grain_858:
XU_858 in out fe_tanh Vc=0.41111741145987635 Qo=2.870840350313312e-13 K=2.62 tau=9.752139286795875e-08 off=-0.1

*Grain_859:
XU_859 in out fe_tanh Vc=0.12063408618438021 Qo=5.831287591493789e-14 K=2.62 tau=8.260593158137339e-08 off=-0.1

*Grain_860:
XU_860 in out fe_tanh Vc=0.32210405628617056 Qo=2.0904917722056366e-13 K=2.62 tau=8.722621849310253e-08 off=-0.1

*Grain_861:
XU_861 in out fe_tanh Vc=0.9039551918298628 Qo=7.995477121793845e-13 K=2.62 tau=1.1239914916696439e-07 off=-0.1

*Grain_862:
XU_862 in out fe_tanh Vc=0.1375624173286063 Qo=6.916767045074323e-14 K=2.62 tau=9.050695434960216e-08 off=-0.1

*Grain_863:
XU_863 in out fe_tanh Vc=0.5916236122359283 Qo=4.608000937975322e-13 K=2.62 tau=9.269546883605072e-08 off=-0.1

*Grain_864:
XU_864 in out fe_tanh Vc=0.42743203281291303 Qo=3.019816796865915e-13 K=2.62 tau=9.952790434371661e-08 off=-0.1

*Grain_865:
XU_865 in out fe_tanh Vc=0.2122643319358916 Qo=1.2156079748059475e-13 K=2.62 tau=1.0972334754423045e-07 off=-0.1

*Grain_866:
XU_866 in out fe_tanh Vc=0.2776355215210951 Qo=1.7233399260475611e-13 K=2.62 tau=9.171581419273263e-08 off=-0.1

*Grain_867:
XU_867 in out fe_tanh Vc=0.4308750790315275 Qo=3.0514776917124303e-13 K=2.62 tau=1.0648009769600064e-07 off=-0.1

*Grain_868:
XU_868 in out fe_tanh Vc=0.22101646210834225 Qo=1.281166045047466e-13 K=2.62 tau=9.517769942816314e-08 off=-0.1

*Grain_869:
XU_869 in out fe_tanh Vc=0.19457619860087896 Qo=1.0856005112146162e-13 K=2.62 tau=9.181654948874255e-08 off=-0.1

*Grain_870:
XU_870 in out fe_tanh Vc=0.4244962493724848 Qo=2.992880833616677e-13 K=2.62 tau=1.0195684996206615e-07 off=-0.1

*Grain_871:
XU_871 in out fe_tanh Vc=0.6151501687180577 Qo=4.847623722959881e-13 K=2.62 tau=1.1198806478801175e-07 off=-0.1

*Grain_872:
XU_872 in out fe_tanh Vc=0.1645485606249502 Qo=8.730431806936831e-14 K=2.62 tau=1.0484525842866132e-07 off=-0.1

*Grain_873:
XU_873 in out fe_tanh Vc=0.5178444966223306 Qo=3.875364754421784e-13 K=2.62 tau=9.724825814930554e-08 off=-0.1

*Grain_874:
XU_874 in out fe_tanh Vc=0.21039861057978837 Qo=1.2017361849111875e-13 K=2.62 tau=1.0390262449294714e-07 off=-0.1

*Grain_875:
XU_875 in out fe_tanh Vc=0.29305167466067444 Qo=1.848761464772846e-13 K=2.62 tau=8.918714403416323e-08 off=-0.1

*Grain_876:
XU_876 in out fe_tanh Vc=0.7681041733465186 Qo=6.469929861411842e-13 K=2.62 tau=1.0229424946750172e-07 off=-0.1

*Grain_877:
XU_877 in out fe_tanh Vc=0.1974723295962157 Qo=1.1066531764411013e-13 K=2.62 tau=8.734894808160631e-08 off=-0.1

*Grain_878:
XU_878 in out fe_tanh Vc=0.16175437558826372 Qo=8.538198734818748e-14 K=2.62 tau=1.1178767332413416e-07 off=-0.1

*Grain_879:
XU_879 in out fe_tanh Vc=1.125529831502031 Qo=1.0632062568122772e-12 K=2.62 tau=8.810890702655473e-08 off=-0.1

*Grain_880:
XU_880 in out fe_tanh Vc=-0.18729420235674 Qo=1.033082595011036e-13 K=2.62 tau=9.406285310440402e-08 off=-0.1

*Grain_881:
XU_881 in out fe_tanh Vc=0.1039860799754973 Qo=4.8075208794411135e-14 K=2.62 tau=9.335028668331591e-08 off=-0.1

*Grain_882:
XU_882 in out fe_tanh Vc=0.7083392367313648 Qo=5.823272311462488e-13 K=2.62 tau=7.993933875855544e-08 off=-0.1

*Grain_883:
XU_883 in out fe_tanh Vc=0.4749566096993875 Qo=3.463406973653688e-13 K=2.62 tau=8.879393457261797e-08 off=-0.1

*Grain_884:
XU_884 in out fe_tanh Vc=0.6623822723799958 Qo=5.336969506034009e-13 K=2.62 tau=8.698022957296285e-08 off=-0.1

*Grain_885:
XU_885 in out fe_tanh Vc=-0.0899727627004634 Qo=3.9828851505048957e-14 K=2.62 tau=1.0602944051887664e-07 off=-0.1

*Grain_886:
XU_886 in out fe_tanh Vc=0.40547615675858795 Qo=2.819735216056334e-13 K=2.62 tau=1.008786473188315e-07 off=-0.1

*Grain_887:
XU_887 in out fe_tanh Vc=0.6750054529443719 Qo=5.469566110924757e-13 K=2.62 tau=1.0528574331566736e-07 off=-0.1

*Grain_888:
XU_888 in out fe_tanh Vc=0.09742934255865504 Qo=4.4172310269743076e-14 K=2.62 tau=8.036757382191194e-08 off=-0.1

*Grain_889:
XU_889 in out fe_tanh Vc=0.47067910078087166 Qo=3.4229125207339153e-13 K=2.62 tau=1.0194878188593857e-07 off=-0.1

*Grain_890:
XU_890 in out fe_tanh Vc=0.332131524694133 Qo=2.1754872350803652e-13 K=2.62 tau=8.602763555794925e-08 off=-0.1

*Grain_891:
XU_891 in out fe_tanh Vc=0.340675211024426 Qo=2.2485166308673295e-13 K=2.62 tau=1.0865524012206506e-07 off=-0.1

*Grain_892:
XU_892 in out fe_tanh Vc=0.5342912919478339 Qo=4.036128040728455e-13 K=2.62 tau=1.0189947465861145e-07 off=-0.1

*Grain_893:
XU_893 in out fe_tanh Vc=0.6076576826556528 Qo=4.771007523917929e-13 K=2.62 tau=9.29635305196394e-08 off=-0.1

*Grain_894:
XU_894 in out fe_tanh Vc=0.4703371014096436 Qo=3.419679621264522e-13 K=2.62 tau=1.0456401528488289e-07 off=-0.1

*Grain_895:
XU_895 in out fe_tanh Vc=0.07554908854315484 Qo=3.173594306840807e-14 K=2.62 tau=9.730564994960743e-08 off=-0.1

*Grain_896:
XU_896 in out fe_tanh Vc=0.797506137775929 Qo=6.793720174998815e-13 K=2.62 tau=9.621853286478218e-08 off=-0.1

*Grain_897:
XU_897 in out fe_tanh Vc=0.16708037744977672 Qo=8.905462771344088e-14 K=2.62 tau=9.802753115703102e-08 off=-0.1

*Grain_898:
XU_898 in out fe_tanh Vc=0.14858132353049885 Qo=7.645517731341251e-14 K=2.62 tau=1.0144220556595431e-07 off=-0.1

*Grain_899:
XU_899 in out fe_tanh Vc=0.49390077757628265 Qo=3.6440559238837326e-13 K=2.62 tau=9.196199195031269e-08 off=-0.1

*Grain_900:
XU_900 in out fe_tanh Vc=0.31556199166523496 Qo=2.0354643736378426e-13 K=2.62 tau=9.143759223976386e-08 off=-0.1

*Grain_901:
XU_901 in out fe_tanh Vc=0.935706480424306 Qo=8.362477049977604e-13 K=2.62 tau=1.0030733448690162e-07 off=-0.1

*Grain_902:
XU_902 in out fe_tanh Vc=0.3916019039103512 Qo=2.694955779610969e-13 K=2.62 tau=1.0229098934582827e-07 off=-0.1

*Grain_903:
XU_903 in out fe_tanh Vc=0.327390610530188 Qo=2.135204598919285e-13 K=2.62 tau=8.392461415182431e-08 off=-0.1

*Grain_904:
XU_904 in out fe_tanh Vc=0.22407002092865372 Qo=1.304224311867345e-13 K=2.62 tau=1.0701061654115687e-07 off=-0.1

*Grain_905:
XU_905 in out fe_tanh Vc=0.7339623995680495 Qo=6.098588996452889e-13 K=2.62 tau=1.036059515906271e-07 off=-0.1

*Grain_906:
XU_906 in out fe_tanh Vc=0.3277285558545808 Qo=2.1380702960828292e-13 K=2.62 tau=1.0345521090190592e-07 off=-0.1

*Grain_907:
XU_907 in out fe_tanh Vc=0.013553582363071748 Qo=3.40035092346308e-15 K=2.62 tau=1.135781281371573e-07 off=-0.1

*Grain_908:
XU_908 in out fe_tanh Vc=0.22009953055876683 Qo=1.2742606193679518e-13 K=2.62 tau=8.920426754147022e-08 off=-0.1

*Grain_909:
XU_909 in out fe_tanh Vc=0.40380461701054954 Qo=2.804633226196333e-13 K=2.62 tau=8.357125426660767e-08 off=-0.1

*Grain_910:
XU_910 in out fe_tanh Vc=0.047012393288290766 Qo=1.7128900210703752e-14 K=2.62 tau=1.0270658367037044e-07 off=-0.1

*Grain_911:
XU_911 in out fe_tanh Vc=0.8201887519858843 Qo=7.045979288861671e-13 K=2.62 tau=1.0620998696882294e-07 off=-0.1

*Grain_912:
XU_912 in out fe_tanh Vc=-0.1820427502791967 Qo=9.955860782353527e-14 K=2.62 tau=1.0330400573882857e-07 off=-0.1

*Grain_913:
XU_913 in out fe_tanh Vc=0.28902561138869703 Qo=1.815810978483189e-13 K=2.62 tau=8.715092291470976e-08 off=-0.1

*Grain_914:
XU_914 in out fe_tanh Vc=0.14481147312990145 Qo=7.394303519566375e-14 K=2.62 tau=1.1952136554674548e-07 off=-0.1

*Grain_915:
XU_915 in out fe_tanh Vc=0.1657477006328489 Qo=8.813231467037244e-14 K=2.62 tau=1.0064233136325628e-07 off=-0.1

*Grain_916:
XU_916 in out fe_tanh Vc=0.6593443145792985 Qo=5.305170619834635e-13 K=2.62 tau=9.488882291742398e-08 off=-0.1

*Grain_917:
XU_917 in out fe_tanh Vc=0.1749707664248677 Qo=9.456023717875036e-14 K=2.62 tau=1.0127760392806984e-07 off=-0.1

*Grain_918:
XU_918 in out fe_tanh Vc=0.2573130081784505 Qo=1.5611825023806085e-13 K=2.62 tau=9.216546715109922e-08 off=-0.1

*Grain_919:
XU_919 in out fe_tanh Vc=-0.007195409150258236 Qo=1.4928822444224896e-15 K=2.62 tau=9.749090716772755e-08 off=-0.1

*Grain_920:
XU_920 in out fe_tanh Vc=-0.06826524523085559 Qo=2.781717108193395e-14 K=2.62 tau=9.587141438147475e-08 off=-0.1

*Grain_921:
XU_921 in out fe_tanh Vc=0.5352603967174361 Qo=4.0456476476457355e-13 K=2.62 tau=1.104483548990806e-07 off=-0.1

*Grain_922:
XU_922 in out fe_tanh Vc=0.2082578000509308 Qo=1.185864504051575e-13 K=2.62 tau=1.2572056483643487e-07 off=-0.1

*Grain_923:
XU_923 in out fe_tanh Vc=0.13394316649190519 Qo=6.681133359540861e-14 K=2.62 tau=9.728006806089813e-08 off=-0.1

*Grain_924:
XU_924 in out fe_tanh Vc=0.5807511970632464 Qo=4.498218611965143e-13 K=2.62 tau=8.854681706513074e-08 off=-0.1

*Grain_925:
XU_925 in out fe_tanh Vc=0.5014554460399276 Qo=3.716682548322763e-13 K=2.62 tau=1.0825953701949966e-07 off=-0.1

*Grain_926:
XU_926 in out fe_tanh Vc=0.9051486162988317 Qo=8.009202418506485e-13 K=2.62 tau=1.072440693278303e-07 off=-0.1

*Grain_927:
XU_927 in out fe_tanh Vc=0.5686949255114193 Qo=4.3772018024650555e-13 K=2.62 tau=8.50397830359055e-08 off=-0.1

*Grain_928:
XU_928 in out fe_tanh Vc=0.4322790736697005 Qo=3.0644101081928464e-13 K=2.62 tau=9.58423976325393e-08 off=-0.1

*Grain_929:
XU_929 in out fe_tanh Vc=0.41930841684406145 Qo=2.945418868675685e-13 K=2.62 tau=9.42033728180075e-08 off=-0.1

*Grain_930:
XU_930 in out fe_tanh Vc=0.32652395468166884 Qo=2.1278596173094406e-13 K=2.62 tau=1.0902839438253644e-07 off=-0.1

*Grain_931:
XU_931 in out fe_tanh Vc=0.4042644375823382 Qo=2.808785736310618e-13 K=2.62 tau=9.54652855078646e-08 off=-0.1

*Grain_932:
XU_932 in out fe_tanh Vc=-0.3087736935644979 Qo=1.9787265960847131e-13 K=2.62 tau=1.0462892453199301e-07 off=-0.1

*Grain_933:
XU_933 in out fe_tanh Vc=0.577772694618771 Qo=4.4682506559384926e-13 K=2.62 tau=8.861391011295783e-08 off=-0.1

*Grain_934:
XU_934 in out fe_tanh Vc=1.0817321271170255 Qo=1.0097388291923662e-12 K=2.62 tau=9.73068040533512e-08 off=-0.1

*Grain_935:
XU_935 in out fe_tanh Vc=0.3577274872604962 Qo=2.3959150524851056e-13 K=2.62 tau=9.146886487596825e-08 off=-0.1

*Grain_936:
XU_936 in out fe_tanh Vc=0.30991933619080714 Qo=1.988276069919328e-13 K=2.62 tau=8.79448404094913e-08 off=-0.1

*Grain_937:
XU_937 in out fe_tanh Vc=0.4372684229852243 Qo=3.1104696026893767e-13 K=2.62 tau=9.662230478827075e-08 off=-0.1

*Grain_938:
XU_938 in out fe_tanh Vc=0.056843871128143986 Qo=2.1925128655601275e-14 K=2.62 tau=9.824338578959204e-08 off=-0.1

*Grain_939:
XU_939 in out fe_tanh Vc=0.37904395834854043 Qo=2.5831514095861665e-13 K=2.62 tau=9.942893728869962e-08 off=-0.1

*Grain_940:
XU_940 in out fe_tanh Vc=0.9256905219284666 Qo=8.246297004211149e-13 K=2.62 tau=1.138296175166806e-07 off=-0.1

*Grain_941:
XU_941 in out fe_tanh Vc=0.23387699371356965 Qo=1.3789139460019655e-13 K=2.62 tau=1.0056546862327694e-07 off=-0.1

*Grain_942:
XU_942 in out fe_tanh Vc=-0.1858938381742351 Qo=1.0230524581397931e-13 K=2.62 tau=8.966229333511031e-08 off=-0.1

*Grain_943:
XU_943 in out fe_tanh Vc=0.6643646219258932 Qo=5.357742753255938e-13 K=2.62 tau=9.424334718453969e-08 off=-0.1

*Grain_944:
XU_944 in out fe_tanh Vc=0.7443654692871686 Qo=6.211199720176372e-13 K=2.62 tau=1.0633342392660877e-07 off=-0.1

*Grain_945:
XU_945 in out fe_tanh Vc=0.5434898354724762 Qo=4.126693980254252e-13 K=2.62 tau=1.0256187192675342e-07 off=-0.1

*Grain_946:
XU_946 in out fe_tanh Vc=0.6625322627203124 Qo=5.338540619003514e-13 K=2.62 tau=1.0386306018820569e-07 off=-0.1

*Grain_947:
XU_947 in out fe_tanh Vc=-0.1038570021044497 Qo=4.799764478969882e-14 K=2.62 tau=1.0284353651737858e-07 off=-0.1

*Grain_948:
XU_948 in out fe_tanh Vc=0.4963197411348312 Qo=3.667274553061338e-13 K=2.62 tau=1.0932991513259022e-07 off=-0.1

*Grain_949:
XU_949 in out fe_tanh Vc=0.3721580452097371 Qo=2.5223133928305217e-13 K=2.62 tau=1.1408095722009696e-07 off=-0.1

*Grain_950:
XU_950 in out fe_tanh Vc=0.4694089555236424 Qo=3.4109094687304363e-13 K=2.62 tau=8.85433906063971e-08 off=-0.1

*Grain_951:
XU_951 in out fe_tanh Vc=0.2466863891978725 Qo=1.4778901514673926e-13 K=2.62 tau=9.231573461321758e-08 off=-0.1

*Grain_952:
XU_952 in out fe_tanh Vc=0.31323069700843503 Qo=2.015937308796463e-13 K=2.62 tau=1.0708836340950891e-07 off=-0.1

*Grain_953:
XU_953 in out fe_tanh Vc=0.3920938854060087 Qo=2.6993580912252413e-13 K=2.62 tau=1.1097923062037043e-07 off=-0.1

*Grain_954:
XU_954 in out fe_tanh Vc=0.1997585518411927 Qo=1.1233378843412871e-13 K=2.62 tau=9.740707219703359e-08 off=-0.1

*Grain_955:
XU_955 in out fe_tanh Vc=1.056842014862 Qo=9.79639982585935e-13 K=2.62 tau=8.898597239686721e-08 off=-0.1

*Grain_956:
XU_956 in out fe_tanh Vc=0.320950423150749 Qo=2.0807636332112802e-13 K=2.62 tau=9.483489787099384e-08 off=-0.1

*Grain_957:
XU_957 in out fe_tanh Vc=0.8497091747616345 Qo=7.377425122349252e-13 K=2.62 tau=1.0249496150298083e-07 off=-0.1

*Grain_958:
XU_958 in out fe_tanh Vc=0.6279882181129973 Qo=4.979552953164794e-13 K=2.62 tau=8.959836713061903e-08 off=-0.1

*Grain_959:
XU_959 in out fe_tanh Vc=0.1757966275357021 Qo=9.514086850155403e-14 K=2.62 tau=8.689477648013266e-08 off=-0.1

*Grain_960:
XU_960 in out fe_tanh Vc=0.6843705343846722 Qo=5.568421529476953e-13 K=2.62 tau=1.0087259429906058e-07 off=-0.1

*Grain_961:
XU_961 in out fe_tanh Vc=0.4434733427266514 Qo=3.167970914877315e-13 K=2.62 tau=1.0471419738861814e-07 off=-0.1

*Grain_962:
XU_962 in out fe_tanh Vc=0.6685741658074313 Qo=5.40191665036682e-13 K=2.62 tau=1.0596216774248935e-07 off=-0.1

*Grain_963:
XU_963 in out fe_tanh Vc=0.6625490415355866 Qo=5.338716379720163e-13 K=2.62 tau=8.851341175280314e-08 off=-0.1

*Grain_964:
XU_964 in out fe_tanh Vc=-0.2572074189962412 Qo=1.5603497268110968e-13 K=2.62 tau=1.0562797440171973e-07 off=-0.1

*Grain_965:
XU_965 in out fe_tanh Vc=0.993349825978183 Qo=9.038290512102649e-13 K=2.62 tau=9.882038191271127e-08 off=-0.1

*Grain_966:
XU_966 in out fe_tanh Vc=0.6149932930379994 Qo=4.846016670277267e-13 K=2.62 tau=9.42051942885738e-08 off=-0.1

*Grain_967:
XU_967 in out fe_tanh Vc=0.25350584386614416 Qo=1.5312206530658725e-13 K=2.62 tau=1.0755624106061544e-07 off=-0.1

*Grain_968:
XU_968 in out fe_tanh Vc=0.246568888863573 Qo=1.4769750939615202e-13 K=2.62 tau=1.1436464041671755e-07 off=-0.1

*Grain_969:
XU_969 in out fe_tanh Vc=0.1593278723654247 Qo=8.372066978325303e-14 K=2.62 tau=7.625131635946763e-08 off=-0.1

*Grain_970:
XU_970 in out fe_tanh Vc=0.49250008758815733 Qo=3.630626858413083e-13 K=2.62 tau=1.1257592102786351e-07 off=-0.1

*Grain_971:
XU_971 in out fe_tanh Vc=0.5651781474559416 Qo=4.3420456037046e-13 K=2.62 tau=8.839545660971644e-08 off=-0.1

*Grain_972:
XU_972 in out fe_tanh Vc=0.6595968507809635 Qo=5.307812292695498e-13 K=2.62 tau=9.47994733923292e-08 off=-0.1

*Grain_973:
XU_973 in out fe_tanh Vc=-0.19242760361104627 Qo=1.0700424160447648e-13 K=2.62 tau=1.0059360645362852e-07 off=-0.1

*Grain_974:
XU_974 in out fe_tanh Vc=0.45430636808077773 Qo=3.268939494375373e-13 K=2.62 tau=9.319492798551566e-08 off=-0.1

*Grain_975:
XU_975 in out fe_tanh Vc=0.2916409669568116 Qo=1.837200262434429e-13 K=2.62 tau=1.0047979175169374e-07 off=-0.1

*Grain_976:
XU_976 in out fe_tanh Vc=0.6456272444927043 Qo=5.162140416461928e-13 K=2.62 tau=1.1154112785011458e-07 off=-0.1

*Grain_977:
XU_977 in out fe_tanh Vc=0.26948717257117616 Qo=1.6578794091438626e-13 K=2.62 tau=1.1113878819814692e-07 off=-0.1

*Grain_978:
XU_978 in out fe_tanh Vc=0.18340672525346263 Qo=1.0052943551908814e-13 K=2.62 tau=1.2149241257307835e-07 off=-0.1

*Grain_979:
XU_979 in out fe_tanh Vc=0.3781396431250376 Qo=2.57514260044201e-13 K=2.62 tau=9.577964235892881e-08 off=-0.1

*Grain_980:
XU_980 in out fe_tanh Vc=0.4717036039685964 Qo=3.4326013042497384e-13 K=2.62 tau=1.1243536835806747e-07 off=-0.1

*Grain_981:
XU_981 in out fe_tanh Vc=0.4769493949096123 Qo=3.4823097853772807e-13 K=2.62 tau=1.1129510098314796e-07 off=-0.1

*Grain_982:
XU_982 in out fe_tanh Vc=0.4966334639516373 Qo=3.6702883396979427e-13 K=2.62 tau=9.233873138881615e-08 off=-0.1

*Grain_983:
XU_983 in out fe_tanh Vc=0.3548546314015615 Qo=2.3709316359097006e-13 K=2.62 tau=1.0537576151411815e-07 off=-0.1

*Grain_984:
XU_984 in out fe_tanh Vc=0.17987765515544404 Qo=9.802205277853658e-14 K=2.62 tau=1.0310820876818245e-07 off=-0.1

*Grain_985:
XU_985 in out fe_tanh Vc=0.7086738629291724 Qo=5.826848824903352e-13 K=2.62 tau=1.0752869972197829e-07 off=-0.1

*Grain_986:
XU_986 in out fe_tanh Vc=0.370899930668698 Qo=2.5112340318527785e-13 K=2.62 tau=1.079949881423852e-07 off=-0.1

*Grain_987:
XU_987 in out fe_tanh Vc=0.6958086491837407 Qo=5.689710640505533e-13 K=2.62 tau=9.96553936961793e-08 off=-0.1

*Grain_988:
XU_988 in out fe_tanh Vc=0.4299669152169913 Qo=3.043119179637322e-13 K=2.62 tau=9.58403099170453e-08 off=-0.1

*Grain_989:
XU_989 in out fe_tanh Vc=0.3939807799070244 Qo=2.7162576137803845e-13 K=2.62 tau=9.282381282316158e-08 off=-0.1

*Grain_990:
XU_990 in out fe_tanh Vc=-0.1935999714408364 Qo=1.0785251728287598e-13 K=2.62 tau=1.116199468282197e-07 off=-0.1

*Grain_991:
XU_991 in out fe_tanh Vc=0.6604010022219258 Qo=5.316226197040235e-13 K=2.62 tau=8.438000691746394e-08 off=-0.1

*Grain_992:
XU_992 in out fe_tanh Vc=0.7540349253925203 Qo=6.316293627934485e-13 K=2.62 tau=1.0653525051848369e-07 off=-0.1

*Grain_993:
XU_993 in out fe_tanh Vc=0.5575670107776701 Qo=4.266184187902257e-13 K=2.62 tau=9.331805539468979e-08 off=-0.1

*Grain_994:
XU_994 in out fe_tanh Vc=0.6253180744899869 Qo=4.952046190317837e-13 K=2.62 tau=1.0972870482880063e-07 off=-0.1

*Grain_995:
XU_995 in out fe_tanh Vc=0.27918188794103893 Qo=1.735828530158153e-13 K=2.62 tau=9.880031732578613e-08 off=-0.1

*Grain_996:
XU_996 in out fe_tanh Vc=0.26377492261949115 Qo=1.6123412535233198e-13 K=2.62 tau=9.26987697035977e-08 off=-0.1

*Grain_997:
XU_997 in out fe_tanh Vc=0.694033225653852 Qo=5.67084466230331e-13 K=2.62 tau=9.90417965074488e-08 off=-0.1

*Grain_998:
XU_998 in out fe_tanh Vc=0.6152108231681065 Qo=4.848245107150163e-13 K=2.62 tau=1.0101174180305553e-07 off=-0.1

*Grain_999:
XU_999 in out fe_tanh Vc=0.19838614255303386 Qo=1.1133152124818536e-13 K=2.62 tau=8.094867529057934e-08 off=-0.1
Rp in out R=50000.0
Cp in out 1.9e-10
.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.ends
