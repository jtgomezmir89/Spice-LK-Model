* Multi-domian SPICE model
V1 in 0 SINE(0 2.1 1k 0 0 0 10)
Rsh 0 N0 0.00000001
B1 Q 0 V=idt(-I(Rsh))

*Grain_0:
XU_0 in N0 fe_tanh Vc=0.9917940605875019 Qo=1.0493510497138771e-07 K=2.62 tau=1.0596447837318364e-08

*Grain_1:
XU_1 in N0 fe_tanh Vc=0.8203206873947178 Qo=7.757001946443028e-08 K=2.62 tau=9.191004048023958e-09

*Grain_2:
XU_2 in N0 fe_tanh Vc=1.0959796774374058 Qo=1.0736293634017652e-07 K=2.62 tau=9.736133245951974e-09

*Grain_3:
XU_3 in N0 fe_tanh Vc=1.0469921631194106 Qo=8.822339812798354e-08 K=2.62 tau=1.1836647919864073e-08

*Grain_4:
XU_4 in N0 fe_tanh Vc=0.9627201753784905 Qo=1.0964906279025674e-07 K=2.62 tau=1.1122584763082123e-08

*Grain_5:
XU_5 in N0 fe_tanh Vc=1.1472767648559812 Qo=9.528055450216515e-08 K=2.62 tau=9.529863222234245e-09

*Grain_6:
XU_6 in N0 fe_tanh Vc=1.0880755043088075 Qo=1.1470775183726527e-07 K=2.62 tau=7.588076000795608e-09

*Grain_7:
XU_7 in N0 fe_tanh Vc=1.0036754963339507 Qo=1.074972642238811e-07 K=2.62 tau=9.545989422965803e-09

*Grain_8:
XU_8 in N0 fe_tanh Vc=1.0616164074075833 Qo=1.060847283076465e-07 K=2.62 tau=9.417946890826759e-09

*Grain_9:
XU_9 in N0 fe_tanh Vc=0.83944176973507 Qo=8.868917943480713e-08 K=2.62 tau=9.502739271743436e-09
Rp in N0 R=1000000000.0Cp in N0 1e-09.tran 0 1.5m 0 1e-8

.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.backanno
.end
