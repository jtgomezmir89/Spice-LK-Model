* Multi-domian SPICE model
V1 in 0 SINE(0 2.1 1k 0 0 0 10)
Rsh 0 N0 0.00000001
B1 Q 0 V=idt(-I(Rsh))

*Grain_0:
XU_0 in N0 fe_tanh Vc=1.0820811594841706 Qo=0.10852541488088509 K=2.62 tau=9.729956249641967e-09

*Grain_1:
XU_1 in N0 fe_tanh Vc=1.0001589273223794 Qo=0.09811023313514114 K=2.62 tau=9.448431255083717e-09

*Grain_2:
XU_2 in N0 fe_tanh Vc=1.0146770863283412 Qo=0.10414155257019891 K=2.62 tau=9.009166804840328e-09

*Grain_3:
XU_3 in N0 fe_tanh Vc=1.0571443323691918 Qo=0.11155168054483452 K=2.62 tau=9.772579678281376e-09

*Grain_4:
XU_4 in N0 fe_tanh Vc=0.9745796814988666 Qo=0.06973685586622871 K=2.62 tau=1.1656655596780314e-08

*Grain_5:
XU_5 in N0 fe_tanh Vc=1.0638487709747901 Qo=0.08880441411722027 K=2.62 tau=9.516948541857998e-09

*Grain_6:
XU_6 in N0 fe_tanh Vc=0.9251567376382758 Qo=0.09214493217005262 K=2.62 tau=8.48454182419285e-09

*Grain_7:
XU_7 in N0 fe_tanh Vc=1.1124685906292286 Qo=0.12368312989104067 K=2.62 tau=1.0253260779798798e-08

*Grain_8:
XU_8 in N0 fe_tanh Vc=1.0339690807537472 Qo=0.10339305598208169 K=2.62 tau=9.470052756198275e-09

*Grain_9:
XU_9 in N0 fe_tanh Vc=0.7295953056419122 Qo=0.09990873084231637 K=2.62 tau=1.007881455660506e-08
.tran 0 1.5m 0 1e-8

.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.backanno
.end
