* Multi-domian SPICE model
.subckt fe_tanh_md in out

*Grain_0:
XU_0 in out fe_tanh Vc=1.0182095080288638 Qo=1.1535894423040818e-07 K=2.62 tau=1.0895113522713204e-08

*Grain_1:
XU_1 in out fe_tanh Vc=0.9421108845199656 Qo=1.0178243509347752e-07 K=2.62 tau=9.370057035967819e-09

*Grain_2:
XU_2 in out fe_tanh Vc=1.0228739469521289 Qo=9.067542653107444e-08 K=2.62 tau=8.580057249636296e-09

*Grain_3:
XU_3 in out fe_tanh Vc=1.0638025883708149 Qo=8.97460424233869e-08 K=2.62 tau=1.0624844702906523e-08

*Grain_4:
XU_4 in out fe_tanh Vc=0.9322003893200547 Qo=9.522004252490078e-08 K=2.62 tau=9.262329478608197e-09

*Grain_5:
XU_5 in out fe_tanh Vc=0.8467065574288073 Qo=1.0458199932441934e-07 K=2.62 tau=1.0154188070604373e-08

*Grain_6:
XU_6 in out fe_tanh Vc=0.8300195156457233 Qo=1.1008109983360041e-07 K=2.62 tau=8.901269312374233e-09

*Grain_7:
XU_7 in out fe_tanh Vc=1.0185167980518053 Qo=9.696253460406616e-08 K=2.62 tau=1.0370826119636214e-08

*Grain_8:
XU_8 in out fe_tanh Vc=1.0190517495549511 Qo=1.0458373164496806e-07 K=2.62 tau=9.587248958996689e-09

*Grain_9:
XU_9 in out fe_tanh Vc=1.1332287252419753 Qo=9.100774378969808e-08 K=2.62 tau=8.641682626924946e-09
Rp in out R=1000000000.0
Cp in out 1e-09
.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.ends
