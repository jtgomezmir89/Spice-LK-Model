* Multi-domian SPICE model
.subckt fe_tanh_md in out

*Grain_0:
XU_0 in out fe_tanh Vc=0.07780821063512039 Qo=2.7434480481591613e-14 K=2.62 tau=9.804763124152627e-08 off=-0.2

*Grain_1:
XU_1 in out fe_tanh Vc=0.35532533717426673 Qo=1.2528454192368148e-13 K=2.62 tau=9.771074966329175e-08 off=-0.2

*Grain_2:
XU_2 in out fe_tanh Vc=0.5314233904330342 Qo=1.8737514348794998e-13 K=2.62 tau=1.174388695545993e-07 off=-0.2

*Grain_3:
XU_3 in out fe_tanh Vc=0.4645101699707024 Qo=1.637821392824827e-13 K=2.62 tau=1.0393505065518789e-07 off=-0.2

*Grain_4:
XU_4 in out fe_tanh Vc=1.1323470127327455 Qo=3.992554483084729e-13 K=2.62 tau=9.581970698504362e-08 off=-0.2

*Grain_5:
XU_5 in out fe_tanh Vc=0.18492934524352816 Qo=6.520443628178085e-14 K=2.62 tau=1.0560977768885068e-07 off=-0.2

*Grain_6:
XU_6 in out fe_tanh Vc=0.31048025613782243 Qo=1.0947256667907404e-13 K=2.62 tau=1.0425079513076926e-07 off=-0.2

*Grain_7:
XU_7 in out fe_tanh Vc=0.36051898953963823 Qo=1.271157773843469e-13 K=2.62 tau=1.0228377471602344e-07 off=-0.2

*Grain_8:
XU_8 in out fe_tanh Vc=0.4391765928062188 Qo=1.5484974612532387e-13 K=2.62 tau=9.013616379809114e-08 off=-0.2

*Grain_9:
XU_9 in out fe_tanh Vc=0.3469030451122352 Qo=1.2231491692781024e-13 K=2.62 tau=9.166048232174367e-08 off=-0.2

*Grain_10:
XU_10 in out fe_tanh Vc=0.5232354572916095 Qo=1.844881513553793e-13 K=2.62 tau=7.548412918751706e-08 off=-0.2

*Grain_11:
XU_11 in out fe_tanh Vc=0.32419929505827927 Qo=1.1430977733354428e-13 K=2.62 tau=1.0323820324713807e-07 off=-0.2

*Grain_12:
XU_12 in out fe_tanh Vc=0.8738937961387272 Qo=3.0812715133086953e-13 K=2.62 tau=1.0551749865726849e-07 off=-0.2

*Grain_13:
XU_13 in out fe_tanh Vc=0.12487232010251392 Qo=4.4028865341843084e-14 K=2.62 tau=1.1646630260416093e-07 off=-0.2

*Grain_14:
XU_14 in out fe_tanh Vc=0.5511527448911273 Qo=1.9433153774733222e-13 K=2.62 tau=9.984080910163287e-08 off=-0.2

*Grain_15:
XU_15 in out fe_tanh Vc=-0.1514045216962821 Qo=5.338388277273277e-14 K=2.62 tau=9.665068554374758e-08 off=-0.2

*Grain_16:
XU_16 in out fe_tanh Vc=0.5454616820815898 Qo=1.923249198044015e-13 K=2.62 tau=1.039712709182433e-07 off=-0.2

*Grain_17:
XU_17 in out fe_tanh Vc=0.6840932983272576 Qo=2.412051901380644e-13 K=2.62 tau=9.796800913153818e-08 off=-0.2

*Grain_18:
XU_18 in out fe_tanh Vc=0.3496643574766144 Qo=1.2328853101745164e-13 K=2.62 tau=1.0505326242721593e-07 off=-0.2

*Grain_19:
XU_19 in out fe_tanh Vc=0.29692287549362206 Qo=1.0469235528969992e-13 K=2.62 tau=8.984538731550499e-08 off=-0.2

*Grain_20:
XU_20 in out fe_tanh Vc=1.2733894773799008 Qo=4.489857622670284e-13 K=2.62 tau=9.673709692950061e-08 off=-0.2

*Grain_21:
XU_21 in out fe_tanh Vc=1.0702328904920926 Qo=3.7735456329476175e-13 K=2.62 tau=9.466823614790931e-08 off=-0.2

*Grain_22:
XU_22 in out fe_tanh Vc=0.5442924836840755 Qo=1.9191267088678868e-13 K=2.62 tau=1.0491061922071995e-07 off=-0.2

*Grain_23:
XU_23 in out fe_tanh Vc=0.28598569075004765 Qo=1.0083600158458442e-13 K=2.62 tau=9.596691571940018e-08 off=-0.2

*Grain_24:
XU_24 in out fe_tanh Vc=0.591328623006003 Qo=2.0849719372343633e-13 K=2.62 tau=1.0741832051514056e-07 off=-0.2

*Grain_25:
XU_25 in out fe_tanh Vc=0.07145892397221287 Qo=2.5195778683880024e-14 K=2.62 tau=1.030452444675879e-07 off=-0.2

*Grain_26:
XU_26 in out fe_tanh Vc=0.5684586580843971 Qo=2.0043344825062527e-13 K=2.62 tau=1.0205386448915763e-07 off=-0.2

*Grain_27:
XU_27 in out fe_tanh Vc=0.43714842210920635 Qo=1.541346312428926e-13 K=2.62 tau=9.450579589239667e-08 off=-0.2

*Grain_28:
XU_28 in out fe_tanh Vc=0.12469030831649203 Qo=4.3964689610898004e-14 K=2.62 tau=9.215030718919846e-08 off=-0.2

*Grain_29:
XU_29 in out fe_tanh Vc=0.5064079749379602 Qo=1.7855493129521844e-13 K=2.62 tau=8.724564630753498e-08 off=-0.2

*Grain_30:
XU_30 in out fe_tanh Vc=0.6913657553658613 Qo=2.437693935691703e-13 K=2.62 tau=9.557732478031654e-08 off=-0.2

*Grain_31:
XU_31 in out fe_tanh Vc=0.506874554627891 Qo=1.7871944312876436e-13 K=2.62 tau=1.0947801486759766e-07 off=-0.2

*Grain_32:
XU_32 in out fe_tanh Vc=0.797620711308139 Qo=2.812339425039973e-13 K=2.62 tau=1.0953734753989458e-07 off=-0.2

*Grain_33:
XU_33 in out fe_tanh Vc=0.8578633491004687 Qo=3.02474958807838e-13 K=2.62 tau=1.0512571996514359e-07 off=-0.2

*Grain_34:
XU_34 in out fe_tanh Vc=0.4663705123720638 Qo=1.6443807940605867e-13 K=2.62 tau=1.0431819523809121e-07 off=-0.2

*Grain_35:
XU_35 in out fe_tanh Vc=0.10064708258121796 Qo=3.5487262848803223e-14 K=2.62 tau=9.1744861108947e-08 off=-0.2

*Grain_36:
XU_36 in out fe_tanh Vc=-0.10038550276876218 Qo=3.539503214203566e-14 K=2.62 tau=9.497154477820546e-08 off=-0.2

*Grain_37:
XU_37 in out fe_tanh Vc=-0.18325007676926514 Qo=6.461234120846571e-14 K=2.62 tau=8.97566424077366e-08 off=-0.2

*Grain_38:
XU_38 in out fe_tanh Vc=1.008130398196274 Qo=3.554577788957794e-13 K=2.62 tau=8.65001002814883e-08 off=-0.2

*Grain_39:
XU_39 in out fe_tanh Vc=0.6137338950412136 Qo=2.163970926327847e-13 K=2.62 tau=1.0902805788556373e-07 off=-0.2

*Grain_40:
XU_40 in out fe_tanh Vc=0.40823901979598565 Qo=1.4394143405942536e-13 K=2.62 tau=1.0426961882209138e-07 off=-0.2

*Grain_41:
XU_41 in out fe_tanh Vc=0.6215757976287541 Qo=2.191620774810459e-13 K=2.62 tau=9.595671954769299e-08 off=-0.2

*Grain_42:
XU_42 in out fe_tanh Vc=0.7314689527545618 Qo=2.579094229700407e-13 K=2.62 tau=1.0096444634073725e-07 off=-0.2

*Grain_43:
XU_43 in out fe_tanh Vc=0.8370602136161993 Qo=2.951399589441927e-13 K=2.62 tau=1.0096646380561798e-07 off=-0.2

*Grain_44:
XU_44 in out fe_tanh Vc=0.16206190330465287 Qo=5.71415803901581e-14 K=2.62 tau=1.08745198869301e-07 off=-0.2

*Grain_45:
XU_45 in out fe_tanh Vc=0.4372452035230428 Qo=1.5416875550545054e-13 K=2.62 tau=9.227371794806026e-08 off=-0.2

*Grain_46:
XU_46 in out fe_tanh Vc=0.16436061756274012 Qo=5.795208651710129e-14 K=2.62 tau=1.1103766242424353e-07 off=-0.2

*Grain_47:
XU_47 in out fe_tanh Vc=0.870064767676688 Qo=3.0677707007661873e-13 K=2.62 tau=1.0068905162667571e-07 off=-0.2

*Grain_48:
XU_48 in out fe_tanh Vc=0.6105620878127682 Qo=2.1527874171853196e-13 K=2.62 tau=1.0773291769543816e-07 off=-0.2

*Grain_49:
XU_49 in out fe_tanh Vc=0.7373931738220174 Qo=2.5999825043332627e-13 K=2.62 tau=1.0503041339648578e-07 off=-0.2

*Grain_50:
XU_50 in out fe_tanh Vc=0.06858511268417516 Qo=2.4182498478026512e-14 K=2.62 tau=1.130795750128404e-07 off=-0.2

*Grain_51:
XU_51 in out fe_tanh Vc=0.5039654755280026 Qo=1.7769372780728558e-13 K=2.62 tau=9.070378494744705e-08 off=-0.2

*Grain_52:
XU_52 in out fe_tanh Vc=0.1854721858423125 Qo=6.539583703101286e-14 K=2.62 tau=1.1803308343927239e-07 off=-0.2

*Grain_53:
XU_53 in out fe_tanh Vc=0.7088666140693556 Qo=2.4994004011910385e-13 K=2.62 tau=9.197284883462544e-08 off=-0.2

*Grain_54:
XU_54 in out fe_tanh Vc=0.3385242125698562 Qo=1.1936061537060845e-13 K=2.62 tau=9.298562483715298e-08 off=-0.2

*Grain_55:
XU_55 in out fe_tanh Vc=0.79227380051477 Qo=2.7934866948974706e-13 K=2.62 tau=1.025963810433958e-07 off=-0.2

*Grain_56:
XU_56 in out fe_tanh Vc=0.7070161417167677 Qo=2.492875800866162e-13 K=2.62 tau=1.0970855216520194e-07 off=-0.2

*Grain_57:
XU_57 in out fe_tanh Vc=-0.013086226765454179 Qo=4.614086737685314e-15 K=2.62 tau=1.0077829044769173e-07 off=-0.2

*Grain_58:
XU_58 in out fe_tanh Vc=0.33910373495613744 Qo=1.1956494979065618e-13 K=2.62 tau=9.375473329240663e-08 off=-0.2

*Grain_59:
XU_59 in out fe_tanh Vc=0.4495820541081736 Qo=1.5851861889158157e-13 K=2.62 tau=8.847799358900804e-08 off=-0.2

*Grain_60:
XU_60 in out fe_tanh Vc=0.2869482622064128 Qo=1.0117539568729197e-13 K=2.62 tau=9.160700510284358e-08 off=-0.2

*Grain_61:
XU_61 in out fe_tanh Vc=1.1457429565787425 Qo=4.039787385239353e-13 K=2.62 tau=1.0629185177004861e-07 off=-0.2

*Grain_62:
XU_62 in out fe_tanh Vc=-0.005319715596429686 Qo=1.8756842305790537e-15 K=2.62 tau=9.299975784499801e-08 off=-0.2

*Grain_63:
XU_63 in out fe_tanh Vc=0.6335623123534395 Qo=2.2338841557020718e-13 K=2.62 tau=1.161744607378158e-07 off=-0.2

*Grain_64:
XU_64 in out fe_tanh Vc=1.128578777709742 Qo=3.979268022781274e-13 K=2.62 tau=1.0414058841889105e-07 off=-0.2

*Grain_65:
XU_65 in out fe_tanh Vc=0.16527948251364571 Qo=5.827607009614867e-14 K=2.62 tau=1.002262457866652e-07 off=-0.2

*Grain_66:
XU_66 in out fe_tanh Vc=0.20473197024407527 Qo=7.218666508035149e-14 K=2.62 tau=9.843458304783698e-08 off=-0.2

*Grain_67:
XU_67 in out fe_tanh Vc=0.4615674928159215 Qo=1.6274457758677622e-13 K=2.62 tau=9.915308933614703e-08 off=-0.2

*Grain_68:
XU_68 in out fe_tanh Vc=0.7274769797956291 Qo=2.565018889407792e-13 K=2.62 tau=1.0230584240764726e-07 off=-0.2

*Grain_69:
XU_69 in out fe_tanh Vc=0.41804492986081737 Qo=1.4739891041162463e-13 K=2.62 tau=7.72526380574373e-08 off=-0.2

*Grain_70:
XU_70 in out fe_tanh Vc=0.9626685252201361 Qo=3.3942832831929383e-13 K=2.62 tau=8.43400258774272e-08 off=-0.2

*Grain_71:
XU_71 in out fe_tanh Vc=0.6766923208199666 Qo=2.385956715369924e-13 K=2.62 tau=1.0004630102274168e-07 off=-0.2

*Grain_72:
XU_72 in out fe_tanh Vc=0.3927019567488002 Qo=1.3846320432724245e-13 K=2.62 tau=1.0425234945380932e-07 off=-0.2

*Grain_73:
XU_73 in out fe_tanh Vc=0.157355305836209 Qo=5.5482076138245014e-14 K=2.62 tau=8.99040442895128e-08 off=-0.2

*Grain_74:
XU_74 in out fe_tanh Vc=0.7903233601762936 Qo=2.7866096163784217e-13 K=2.62 tau=9.637966528479385e-08 off=-0.2

*Grain_75:
XU_75 in out fe_tanh Vc=0.9937352227191192 Qo=3.5038216852724043e-13 K=2.62 tau=9.752763129207661e-08 off=-0.2

*Grain_76:
XU_76 in out fe_tanh Vc=0.154909423944543 Qo=5.4619680017456936e-14 K=2.62 tau=9.508251584138256e-08 off=-0.2

*Grain_77:
XU_77 in out fe_tanh Vc=0.40890245835297323 Qo=1.4417535657215047e-13 K=2.62 tau=1.0787823924881604e-07 off=-0.2

*Grain_78:
XU_78 in out fe_tanh Vc=0.2723074666630424 Qo=9.60131818760381e-14 K=2.62 tau=9.83738895416374e-08 off=-0.2

*Grain_79:
XU_79 in out fe_tanh Vc=-0.14152526498763046 Qo=4.990054504868285e-14 K=2.62 tau=9.562457859868135e-08 off=-0.2

*Grain_80:
XU_80 in out fe_tanh Vc=0.8768642055091864 Qo=3.091744911582607e-13 K=2.62 tau=8.936691167929023e-08 off=-0.2

*Grain_81:
XU_81 in out fe_tanh Vc=0.5940061943299828 Qo=2.0944128146978323e-13 K=2.62 tau=8.803938482227676e-08 off=-0.2

*Grain_82:
XU_82 in out fe_tanh Vc=0.7307161391756278 Qo=2.576439876224218e-13 K=2.62 tau=1.0341290241517017e-07 off=-0.2

*Grain_83:
XU_83 in out fe_tanh Vc=0.09181086971337193 Qo=3.2371693071843326e-14 K=2.62 tau=9.572448951029819e-08 off=-0.2

*Grain_84:
XU_84 in out fe_tanh Vc=0.13588087530295828 Qo=4.791038363293194e-14 K=2.62 tau=9.86089050618082e-08 off=-0.2

*Grain_85:
XU_85 in out fe_tanh Vc=0.16240609736079042 Qo=5.72629401417564e-14 K=2.62 tau=9.837871326322018e-08 off=-0.2

*Grain_86:
XU_86 in out fe_tanh Vc=1.0014454778825224 Qo=3.5310073566895797e-13 K=2.62 tau=9.776049417427542e-08 off=-0.2

*Grain_87:
XU_87 in out fe_tanh Vc=0.5358964266710781 Qo=1.8895229613500847e-13 K=2.62 tau=9.542285527729491e-08 off=-0.2

*Grain_88:
XU_88 in out fe_tanh Vc=0.3885534192751014 Qo=1.3700046704771464e-13 K=2.62 tau=1.2017824824252404e-07 off=-0.2

*Grain_89:
XU_89 in out fe_tanh Vc=0.3883893713673554 Qo=1.3694262521988741e-13 K=2.62 tau=9.95323301441307e-08 off=-0.2

*Grain_90:
XU_90 in out fe_tanh Vc=0.7047440776387799 Qo=2.484864705752718e-13 K=2.62 tau=8.468998745438465e-08 off=-0.2

*Grain_91:
XU_91 in out fe_tanh Vc=0.751354722050124 Qo=2.6492096770481044e-13 K=2.62 tau=9.115578663954891e-08 off=-0.2

*Grain_92:
XU_92 in out fe_tanh Vc=0.2599829937369377 Qo=9.166768274198517e-14 K=2.62 tau=1.1159280755583954e-07 off=-0.2

*Grain_93:
XU_93 in out fe_tanh Vc=-0.28528692673896877 Qo=1.0058962363209454e-13 K=2.62 tau=9.875279516703663e-08 off=-0.2

*Grain_94:
XU_94 in out fe_tanh Vc=0.5089339531578689 Qo=1.7944556866633066e-13 K=2.62 tau=8.272497582041194e-08 off=-0.2

*Grain_95:
XU_95 in out fe_tanh Vc=0.8426519949295326 Qo=2.971115711178407e-13 K=2.62 tau=1.0123165955693959e-07 off=-0.2

*Grain_96:
XU_96 in out fe_tanh Vc=0.6184699666734316 Qo=2.1806698921173078e-13 K=2.62 tau=1.234814697618337e-07 off=-0.2

*Grain_97:
XU_97 in out fe_tanh Vc=1.1329690591158004 Qo=3.994747763101743e-13 K=2.62 tau=1.1737379433208077e-07 off=-0.2

*Grain_98:
XU_98 in out fe_tanh Vc=1.0753974450722856 Qo=3.791755391361271e-13 K=2.62 tau=1.1156275655627755e-07 off=-0.2

*Grain_99:
XU_99 in out fe_tanh Vc=0.18684375913109935 Qo=6.587944152870209e-14 K=2.62 tau=7.409569783137805e-08 off=-0.2

*Grain_100:
XU_100 in out fe_tanh Vc=0.4472527795702959 Qo=1.5769733748279375e-13 K=2.62 tau=9.541127793443773e-08 off=-0.2

*Grain_101:
XU_101 in out fe_tanh Vc=0.19752287176943062 Qo=6.964480131330017e-14 K=2.62 tau=1.0140298348337182e-07 off=-0.2

*Grain_102:
XU_102 in out fe_tanh Vc=0.26370843676567407 Qo=9.298124069715316e-14 K=2.62 tau=1.0973901833018787e-07 off=-0.2

*Grain_103:
XU_103 in out fe_tanh Vc=0.0030652796272299665 Qo=1.0807902330284813e-15 K=2.62 tau=8.32744524192486e-08 off=-0.2

*Grain_104:
XU_104 in out fe_tanh Vc=0.9166765440144701 Qo=3.232119663133148e-13 K=2.62 tau=9.271298442502582e-08 off=-0.2

*Grain_105:
XU_105 in out fe_tanh Vc=1.0422160901786959 Qo=3.67476089608238e-13 K=2.62 tau=9.051074170946301e-08 off=-0.2

*Grain_106:
XU_106 in out fe_tanh Vc=0.7620757192084293 Qo=2.6870109559725125e-13 K=2.62 tau=8.295991880307153e-08 off=-0.2

*Grain_107:
XU_107 in out fe_tanh Vc=0.6224481865969188 Qo=2.194696740434666e-13 K=2.62 tau=1.0989729191986353e-07 off=-0.2

*Grain_108:
XU_108 in out fe_tanh Vc=-0.23508784431134094 Qo=8.288987529174469e-14 K=2.62 tau=9.473284543606496e-08 off=-0.2

*Grain_109:
XU_109 in out fe_tanh Vc=0.6795852708951376 Qo=2.396156999083386e-13 K=2.62 tau=1.2106234532747563e-07 off=-0.2

*Grain_110:
XU_110 in out fe_tanh Vc=0.4361308678243095 Qo=1.5377585068567253e-13 K=2.62 tau=9.634339981477336e-08 off=-0.2

*Grain_111:
XU_111 in out fe_tanh Vc=0.6396679440724778 Qo=2.2554120680980082e-13 K=2.62 tau=1.0339216398239941e-07 off=-0.2

*Grain_112:
XU_112 in out fe_tanh Vc=0.27664148378031894 Qo=9.754131762212784e-14 K=2.62 tau=1.1566780656706332e-07 off=-0.2

*Grain_113:
XU_113 in out fe_tanh Vc=1.1685988297541925 Qo=4.120375153728478e-13 K=2.62 tau=1.0063993826082014e-07 off=-0.2

*Grain_114:
XU_114 in out fe_tanh Vc=-0.2181505810839472 Qo=7.691794747550754e-14 K=2.62 tau=8.63594796399289e-08 off=-0.2

*Grain_115:
XU_115 in out fe_tanh Vc=-0.3048283868164989 Qo=1.0747976801021005e-13 K=2.62 tau=9.81145323322743e-08 off=-0.2

*Grain_116:
XU_116 in out fe_tanh Vc=0.3438205024565624 Qo=1.2122803990505866e-13 K=2.62 tau=1.0113878443844883e-07 off=-0.2

*Grain_117:
XU_117 in out fe_tanh Vc=0.3108693895347555 Qo=1.0960977164106654e-13 K=2.62 tau=7.39226988053554e-08 off=-0.2

*Grain_118:
XU_118 in out fe_tanh Vc=0.5183505577074803 Qo=1.8276577936916582e-13 K=2.62 tau=1.1187867736211144e-07 off=-0.2

*Grain_119:
XU_119 in out fe_tanh Vc=0.4986048316732179 Qo=1.7580361263817418e-13 K=2.62 tau=1.0216418798999235e-07 off=-0.2

*Grain_120:
XU_120 in out fe_tanh Vc=-0.34508831566777615 Qo=1.2167505952565443e-13 K=2.62 tau=1.0824482015052401e-07 off=-0.2

*Grain_121:
XU_121 in out fe_tanh Vc=-0.004455668264814916 Qo=1.571028854740644e-15 K=2.62 tau=1.0676234035099276e-07 off=-0.2

*Grain_122:
XU_122 in out fe_tanh Vc=0.31750454723774557 Qo=1.1194926901556083e-13 K=2.62 tau=1.0435538517973437e-07 off=-0.2

*Grain_123:
XU_123 in out fe_tanh Vc=0.37406927543056495 Qo=1.318934872270511e-13 K=2.62 tau=1.0072103665268014e-07 off=-0.2

*Grain_124:
XU_124 in out fe_tanh Vc=0.6315099267959101 Qo=2.226647627441219e-13 K=2.62 tau=8.821196977466854e-08 off=-0.2

*Grain_125:
XU_125 in out fe_tanh Vc=0.35414178980563066 Qo=1.2486723368694342e-13 K=2.62 tau=9.966477062622218e-08 off=-0.2

*Grain_126:
XU_126 in out fe_tanh Vc=0.4142816514477981 Qo=1.4607201203771227e-13 K=2.62 tau=9.20258789123082e-08 off=-0.2

*Grain_127:
XU_127 in out fe_tanh Vc=0.3654144980142052 Qo=1.2884188997062392e-13 K=2.62 tau=1.0553456513045044e-07 off=-0.2

*Grain_128:
XU_128 in out fe_tanh Vc=0.13906557566256705 Qo=4.9033280550136825e-14 K=2.62 tau=1.0032911398551144e-07 off=-0.2

*Grain_129:
XU_129 in out fe_tanh Vc=0.7910289180613337 Qo=2.7890973504964235e-13 K=2.62 tau=1.0189839045593642e-07 off=-0.2

*Grain_130:
XU_130 in out fe_tanh Vc=0.609335265147395 Qo=2.1484617499847989e-13 K=2.62 tau=8.576156085107479e-08 off=-0.2

*Grain_131:
XU_131 in out fe_tanh Vc=0.1485158833299296 Qo=5.236537467142573e-14 K=2.62 tau=8.502433716500449e-08 off=-0.2

*Grain_132:
XU_132 in out fe_tanh Vc=0.5919237530856629 Qo=2.0870703127684064e-13 K=2.62 tau=1.0217396258839339e-07 off=-0.2

*Grain_133:
XU_133 in out fe_tanh Vc=0.5588268136601166 Qo=1.9703734588941278e-13 K=2.62 tau=1.1259561273860159e-07 off=-0.2

*Grain_134:
XU_134 in out fe_tanh Vc=1.1108898375288991 Qo=3.9168983987827066e-13 K=2.62 tau=1.0208650020838426e-07 off=-0.2

*Grain_135:
XU_135 in out fe_tanh Vc=0.6444897647202088 Qo=2.272413377261414e-13 K=2.62 tau=1.0610444338395787e-07 off=-0.2

*Grain_136:
XU_136 in out fe_tanh Vc=0.38133113414744385 Qo=1.3445395378452728e-13 K=2.62 tau=1.1520278555235851e-07 off=-0.2

*Grain_137:
XU_137 in out fe_tanh Vc=0.49801941947794803 Qo=1.7559720152405496e-13 K=2.62 tau=1.1447421728048e-07 off=-0.2

*Grain_138:
XU_138 in out fe_tanh Vc=0.8939233614629779 Qo=3.1518939726169795e-13 K=2.62 tau=9.174448813748025e-08 off=-0.2

*Grain_139:
XU_139 in out fe_tanh Vc=0.7501414534822956 Qo=2.644931800385562e-13 K=2.62 tau=8.692631028398895e-08 off=-0.2

*Grain_140:
XU_140 in out fe_tanh Vc=0.11796598729581786 Qo=4.1593754046542884e-14 K=2.62 tau=9.645598075675096e-08 off=-0.2

*Grain_141:
XU_141 in out fe_tanh Vc=0.3178129718990282 Qo=1.1205801679784411e-13 K=2.62 tau=9.570160822025567e-08 off=-0.2

*Grain_142:
XU_142 in out fe_tanh Vc=0.32528928836904747 Qo=1.1469409924462853e-13 K=2.62 tau=1.0366239629389836e-07 off=-0.2

*Grain_143:
XU_143 in out fe_tanh Vc=0.7168900419497365 Qo=2.527690291651572e-13 K=2.62 tau=1.0344855103245579e-07 off=-0.2

*Grain_144:
XU_144 in out fe_tanh Vc=0.7591867325053137 Qo=2.676824646755111e-13 K=2.62 tau=9.379365595842745e-08 off=-0.2

*Grain_145:
XU_145 in out fe_tanh Vc=0.8100771440404263 Qo=2.8562596948771446e-13 K=2.62 tau=8.865049569009827e-08 off=-0.2

*Grain_146:
XU_146 in out fe_tanh Vc=0.2736922675064798 Qo=9.650145029141568e-14 K=2.62 tau=9.599260173356238e-08 off=-0.2

*Grain_147:
XU_147 in out fe_tanh Vc=0.2426283465158841 Qo=8.554858905554075e-14 K=2.62 tau=9.956199805896202e-08 off=-0.2

*Grain_148:
XU_148 in out fe_tanh Vc=-0.11549007675483963 Qo=4.0720770092070925e-14 K=2.62 tau=8.438433853600005e-08 off=-0.2

*Grain_149:
XU_149 in out fe_tanh Vc=-0.010032060985238012 Qo=3.5372151479013783e-15 K=2.62 tau=1.0502017795665994e-07 off=-0.2

*Grain_150:
XU_150 in out fe_tanh Vc=-0.05165450288995094 Qo=1.821291660293023e-14 K=2.62 tau=9.400493677524426e-08 off=-0.2

*Grain_151:
XU_151 in out fe_tanh Vc=0.8551516015057042 Qo=3.015188208135016e-13 K=2.62 tau=9.681315251947464e-08 off=-0.2

*Grain_152:
XU_152 in out fe_tanh Vc=0.5332218416313317 Qo=1.8800926132582396e-13 K=2.62 tau=7.967287930848973e-08 off=-0.2

*Grain_153:
XU_153 in out fe_tanh Vc=-0.1689112607798549 Qo=5.955660269218824e-14 K=2.62 tau=8.982576877886718e-08 off=-0.2

*Grain_154:
XU_154 in out fe_tanh Vc=0.1773090635751095 Qo=6.251759299120788e-14 K=2.62 tau=1.1505620711980086e-07 off=-0.2

*Grain_155:
XU_155 in out fe_tanh Vc=0.5145370731037581 Qo=1.814211787405987e-13 K=2.62 tau=1.1351443129889518e-07 off=-0.2

*Grain_156:
XU_156 in out fe_tanh Vc=0.10803401509161775 Qo=3.809182930935005e-14 K=2.62 tau=1.215256149345005e-07 off=-0.2

*Grain_157:
XU_157 in out fe_tanh Vc=0.48815839681512885 Qo=1.7212029296179154e-13 K=2.62 tau=1.0992559516936093e-07 off=-0.2

*Grain_158:
XU_158 in out fe_tanh Vc=0.6059221502159151 Qo=2.1364274114227387e-13 K=2.62 tau=8.669607964290323e-08 off=-0.2

*Grain_159:
XU_159 in out fe_tanh Vc=0.8572778037384656 Qo=3.0226850074031744e-13 K=2.62 tau=1.0501388980861631e-07 off=-0.2

*Grain_160:
XU_160 in out fe_tanh Vc=0.6179550956255035 Qo=2.178854502764485e-13 K=2.62 tau=8.728927656659247e-08 off=-0.2

*Grain_161:
XU_161 in out fe_tanh Vc=0.23691088442915428 Qo=8.353266296313645e-14 K=2.62 tau=9.161859746265269e-08 off=-0.2

*Grain_162:
XU_162 in out fe_tanh Vc=0.4980995748033641 Qo=1.756254635762558e-13 K=2.62 tau=9.127045258192862e-08 off=-0.2

*Grain_163:
XU_163 in out fe_tanh Vc=0.09235957377589221 Qo=3.2565161226045916e-14 K=2.62 tau=9.856030601645953e-08 off=-0.2

*Grain_164:
XU_164 in out fe_tanh Vc=0.009132936532871394 Qo=3.220191892416825e-15 K=2.62 tau=1.0538247691537314e-07 off=-0.2

*Grain_165:
XU_165 in out fe_tanh Vc=0.48683137997341586 Qo=1.7165239866958836e-13 K=2.62 tau=1.0319186364475785e-07 off=-0.2

*Grain_166:
XU_166 in out fe_tanh Vc=0.5338678737175532 Qo=1.8823704647234326e-13 K=2.62 tau=1.0608180803765365e-07 off=-0.2

*Grain_167:
XU_167 in out fe_tanh Vc=0.4182310292306856 Qo=1.4746452738814436e-13 K=2.62 tau=1.0057949508895772e-07 off=-0.2

*Grain_168:
XU_168 in out fe_tanh Vc=0.5798219687469053 Qo=2.044400501507611e-13 K=2.62 tau=1.153540405746669e-07 off=-0.2

*Grain_169:
XU_169 in out fe_tanh Vc=0.9622940880605744 Qo=3.392963051194062e-13 K=2.62 tau=9.353354853196293e-08 off=-0.2

*Grain_170:
XU_170 in out fe_tanh Vc=0.01643566970629995 Qo=5.795070418389077e-15 K=2.62 tau=1.0163640576145758e-07 off=-0.2

*Grain_171:
XU_171 in out fe_tanh Vc=0.7239765363069319 Qo=2.5526766381487416e-13 K=2.62 tau=1.1562382197138418e-07 off=-0.2

*Grain_172:
XU_172 in out fe_tanh Vc=0.7264046430059918 Qo=2.561237925614272e-13 K=2.62 tau=9.188943736457602e-08 off=-0.2

*Grain_173:
XU_173 in out fe_tanh Vc=0.18593690281290792 Qo=6.555969208634954e-14 K=2.62 tau=9.982483067134278e-08 off=-0.2

*Grain_174:
XU_174 in out fe_tanh Vc=0.18245859189115055 Qo=6.433327070597161e-14 K=2.62 tau=8.370759473260427e-08 off=-0.2

*Grain_175:
XU_175 in out fe_tanh Vc=0.35403889066812855 Qo=1.2483095236963345e-13 K=2.62 tau=1.102143019495946e-07 off=-0.2

*Grain_176:
XU_176 in out fe_tanh Vc=0.567746096927934 Qo=2.0018220554783905e-13 K=2.62 tau=1.192442290490988e-07 off=-0.2

*Grain_177:
XU_177 in out fe_tanh Vc=1.3109115345044866 Qo=4.622157046524272e-13 K=2.62 tau=7.973998487853772e-08 off=-0.2

*Grain_178:
XU_178 in out fe_tanh Vc=0.2623828597087265 Qo=9.251385406020537e-14 K=2.62 tau=1.152829843113132e-07 off=-0.2

*Grain_179:
XU_179 in out fe_tanh Vc=0.12288189151657547 Qo=4.332705799085534e-14 K=2.62 tau=1.1107078234506429e-07 off=-0.2

*Grain_180:
XU_180 in out fe_tanh Vc=0.3827785460285788 Qo=1.3496429829287274e-13 K=2.62 tau=1.1462439535563688e-07 off=-0.2

*Grain_181:
XU_181 in out fe_tanh Vc=0.3866260737879802 Qo=1.3632090223423155e-13 K=2.62 tau=1.0238255390768587e-07 off=-0.2

*Grain_182:
XU_182 in out fe_tanh Vc=0.20556769661005747 Qo=7.24813347365271e-14 K=2.62 tau=1.0551326829219802e-07 off=-0.2

*Grain_183:
XU_183 in out fe_tanh Vc=0.8838583346907256 Qo=3.1164055867157855e-13 K=2.62 tau=8.915972696651846e-08 off=-0.2

*Grain_184:
XU_184 in out fe_tanh Vc=0.18483826168129075 Qo=6.517232103083241e-14 K=2.62 tau=7.902282588321828e-08 off=-0.2

*Grain_185:
XU_185 in out fe_tanh Vc=0.6311496122101968 Qo=2.2253771903770204e-13 K=2.62 tau=9.596221979150287e-08 off=-0.2

*Grain_186:
XU_186 in out fe_tanh Vc=0.4695713567019867 Qo=1.6556666854308024e-13 K=2.62 tau=1.0820345417268831e-07 off=-0.2

*Grain_187:
XU_187 in out fe_tanh Vc=0.33425288562055977 Qo=1.1785458361811784e-13 K=2.62 tau=1.0577574524705719e-07 off=-0.2

*Grain_188:
XU_188 in out fe_tanh Vc=0.5495310128596542 Qo=1.937597295101211e-13 K=2.62 tau=1.0355182416838313e-07 off=-0.2

*Grain_189:
XU_189 in out fe_tanh Vc=0.47887353298612945 Qo=1.6884653286100412e-13 K=2.62 tau=1.0577964805772853e-07 off=-0.2

*Grain_190:
XU_190 in out fe_tanh Vc=0.9216423056993726 Qo=3.249628495544107e-13 K=2.62 tau=1.0901512092305218e-07 off=-0.2

*Grain_191:
XU_191 in out fe_tanh Vc=0.4433316345901645 Qo=1.563147767665812e-13 K=2.62 tau=9.198878384763537e-08 off=-0.2

*Grain_192:
XU_192 in out fe_tanh Vc=0.8058810714954798 Qo=2.841464717664069e-13 K=2.62 tau=7.106945990235395e-08 off=-0.2

*Grain_193:
XU_193 in out fe_tanh Vc=0.3509534928197412 Qo=1.237430686314188e-13 K=2.62 tau=7.950129547202375e-08 off=-0.2

*Grain_194:
XU_194 in out fe_tanh Vc=1.0067078248214478 Qo=3.549561922230269e-13 K=2.62 tau=9.021685903798106e-08 off=-0.2

*Grain_195:
XU_195 in out fe_tanh Vc=0.6197296077389497 Qo=2.1851112740670647e-13 K=2.62 tau=1.0921604046334205e-07 off=-0.2

*Grain_196:
XU_196 in out fe_tanh Vc=0.08999420702075761 Qo=3.173115402364592e-14 K=2.62 tau=7.709830581837974e-08 off=-0.2

*Grain_197:
XU_197 in out fe_tanh Vc=1.1397609626002885 Qo=4.018695408479664e-13 K=2.62 tau=1.0475288475077843e-07 off=-0.2

*Grain_198:
XU_198 in out fe_tanh Vc=0.24826777189618823 Qo=8.753700010188747e-14 K=2.62 tau=1.059272020835464e-07 off=-0.2

*Grain_199:
XU_199 in out fe_tanh Vc=0.256925847156959 Qo=9.058976014881434e-14 K=2.62 tau=1.1399199746932684e-07 off=-0.2

*Grain_200:
XU_200 in out fe_tanh Vc=0.6760117059879575 Qo=2.383556928230261e-13 K=2.62 tau=1.032885717926576e-07 off=-0.2

*Grain_201:
XU_201 in out fe_tanh Vc=0.7359571966487488 Qo=2.5949193770089765e-13 K=2.62 tau=1.0426668164550712e-07 off=-0.2

*Grain_202:
XU_202 in out fe_tanh Vc=0.5644502874248298 Qo=1.9902013253850109e-13 K=2.62 tau=9.967895468997303e-08 off=-0.2

*Grain_203:
XU_203 in out fe_tanh Vc=0.7664229942511654 Qo=2.7023390596950553e-13 K=2.62 tau=9.203487838401884e-08 off=-0.2

*Grain_204:
XU_204 in out fe_tanh Vc=0.25713326372568723 Qo=9.0662893379355e-14 K=2.62 tau=1.0115969954102201e-07 off=-0.2

*Grain_205:
XU_205 in out fe_tanh Vc=0.09369913315667922 Qo=3.3037477905560277e-14 K=2.62 tau=1.0103942919850472e-07 off=-0.2

*Grain_206:
XU_206 in out fe_tanh Vc=0.35614590603378105 Qo=1.255738671783865e-13 K=2.62 tau=1.1245045470175065e-07 off=-0.2

*Grain_207:
XU_207 in out fe_tanh Vc=0.31494977193170104 Qo=1.1104847804894664e-13 K=2.62 tau=1.1798787934363464e-07 off=-0.2

*Grain_208:
XU_208 in out fe_tanh Vc=0.5023835997581145 Qo=1.771359725321153e-13 K=2.62 tau=9.967727790196817e-08 off=-0.2

*Grain_209:
XU_209 in out fe_tanh Vc=0.23587400743220577 Qo=8.316706939013946e-14 K=2.62 tau=8.293975320391047e-08 off=-0.2

*Grain_210:
XU_210 in out fe_tanh Vc=0.5648006318586446 Qo=1.991436608583644e-13 K=2.62 tau=1.0165240439279178e-07 off=-0.2

*Grain_211:
XU_211 in out fe_tanh Vc=0.18696631694937899 Qo=6.592265432136258e-14 K=2.62 tau=9.837072073418958e-08 off=-0.2

*Grain_212:
XU_212 in out fe_tanh Vc=0.2573076868019383 Qo=9.072439339897874e-14 K=2.62 tau=1.0489078005654931e-07 off=-0.2

*Grain_213:
XU_213 in out fe_tanh Vc=0.734734109025871 Qo=2.59060687923487e-13 K=2.62 tau=1.1699518932358555e-07 off=-0.2

*Grain_214:
XU_214 in out fe_tanh Vc=0.28310666323868994 Qo=9.982088218495312e-14 K=2.62 tau=9.584815130497923e-08 off=-0.2

*Grain_215:
XU_215 in out fe_tanh Vc=0.17331355393907777 Qo=6.110881196117289e-14 K=2.62 tau=1.0109423737596254e-07 off=-0.2

*Grain_216:
XU_216 in out fe_tanh Vc=0.20275213468131228 Qo=7.148859273477224e-14 K=2.62 tau=1.0935168674091519e-07 off=-0.2

*Grain_217:
XU_217 in out fe_tanh Vc=0.9731433337175883 Qo=3.431216522876264e-13 K=2.62 tau=1.0725914730788655e-07 off=-0.2

*Grain_218:
XU_218 in out fe_tanh Vc=0.054861706462336624 Qo=1.9343747952075674e-14 K=2.62 tau=1.0860069844416413e-07 off=-0.2

*Grain_219:
XU_219 in out fe_tanh Vc=0.28995066542116643 Qo=1.0223401625857456e-13 K=2.62 tau=9.597194632931487e-08 off=-0.2

*Grain_220:
XU_220 in out fe_tanh Vc=0.44944149685687423 Qo=1.58469059659518e-13 K=2.62 tau=1.0044212887252138e-07 off=-0.2

*Grain_221:
XU_221 in out fe_tanh Vc=0.35139885300660745 Qo=1.239000986576092e-13 K=2.62 tau=1.0280804955845925e-07 off=-0.2

*Grain_222:
XU_222 in out fe_tanh Vc=0.5653488722155737 Qo=1.99336965514115e-13 K=2.62 tau=1.0864676193714796e-07 off=-0.2

*Grain_223:
XU_223 in out fe_tanh Vc=0.36492045029170234 Qo=1.2866769315399822e-13 K=2.62 tau=8.486571388157162e-08 off=-0.2

*Grain_224:
XU_224 in out fe_tanh Vc=0.330726582212965 Qo=1.1661124051565916e-13 K=2.62 tau=1.0059366654785825e-07 off=-0.2

*Grain_225:
XU_225 in out fe_tanh Vc=0.7702224085289403 Qo=2.7157354552674836e-13 K=2.62 tau=1.247564172839839e-07 off=-0.2

*Grain_226:
XU_226 in out fe_tanh Vc=0.1390007432329587 Qo=4.9010421214211396e-14 K=2.62 tau=1.0376004915120682e-07 off=-0.2

*Grain_227:
XU_227 in out fe_tanh Vc=0.42565832329747755 Qo=1.5008332497317033e-13 K=2.62 tau=1.0563537555357461e-07 off=-0.2

*Grain_228:
XU_228 in out fe_tanh Vc=0.7246404315970663 Qo=2.555017473676296e-13 K=2.62 tau=1.0406861136109312e-07 off=-0.2

*Grain_229:
XU_229 in out fe_tanh Vc=0.47934239452770105 Qo=1.6901184925506874e-13 K=2.62 tau=1.156723766976775e-07 off=-0.2

*Grain_230:
XU_230 in out fe_tanh Vc=0.40026622013302504 Qo=1.4113029607087992e-13 K=2.62 tau=1.0446670066236906e-07 off=-0.2

*Grain_231:
XU_231 in out fe_tanh Vc=0.7926557509695882 Qo=2.7948334181047144e-13 K=2.62 tau=1.0142039964635979e-07 off=-0.2

*Grain_232:
XU_232 in out fe_tanh Vc=0.6441744786625684 Qo=2.271301706767536e-13 K=2.62 tau=8.20565455142899e-08 off=-0.2

*Grain_233:
XU_233 in out fe_tanh Vc=0.2281260045379838 Qo=8.043519273550651e-14 K=2.62 tau=1.1109390198585187e-07 off=-0.2

*Grain_234:
XU_234 in out fe_tanh Vc=0.1345073983401639 Qo=4.742610791678162e-14 K=2.62 tau=1.2115214341141572e-07 off=-0.2

*Grain_235:
XU_235 in out fe_tanh Vc=0.05441314101346417 Qo=1.9185587779115047e-14 K=2.62 tau=1.1161214975976381e-07 off=-0.2

*Grain_236:
XU_236 in out fe_tanh Vc=1.0343396453069011 Qo=3.6469892545890534e-13 K=2.62 tau=9.508259651687509e-08 off=-0.2

*Grain_237:
XU_237 in out fe_tanh Vc=1.0838521312363558 Qo=3.821565860031973e-13 K=2.62 tau=1.09247034681976e-07 off=-0.2

*Grain_238:
XU_238 in out fe_tanh Vc=0.3772521735641783 Qo=1.3301574869545832e-13 K=2.62 tau=1.1337881373665854e-07 off=-0.2

*Grain_239:
XU_239 in out fe_tanh Vc=0.5128598458144668 Qo=1.8082980337088308e-13 K=2.62 tau=9.81275491543143e-08 off=-0.2

*Grain_240:
XU_240 in out fe_tanh Vc=0.4094066101249425 Qo=1.443531159864199e-13 K=2.62 tau=9.37255898189315e-08 off=-0.2

*Grain_241:
XU_241 in out fe_tanh Vc=0.29959467601168605 Qo=1.0563440830139644e-13 K=2.62 tau=9.442431396705272e-08 off=-0.2

*Grain_242:
XU_242 in out fe_tanh Vc=0.5950102402811205 Qo=2.097952991091077e-13 K=2.62 tau=1.0806320238453744e-07 off=-0.2

*Grain_243:
XU_243 in out fe_tanh Vc=0.5874946808043999 Qo=2.0714537992847993e-13 K=2.62 tau=1.0026351310382967e-07 off=-0.2

*Grain_244:
XU_244 in out fe_tanh Vc=0.14641184056948936 Qo=5.1623507976734294e-14 K=2.62 tau=9.879934140785624e-08 off=-0.2

*Grain_245:
XU_245 in out fe_tanh Vc=0.7976611969213091 Qo=2.812482173697889e-13 K=2.62 tau=9.611323773807702e-08 off=-0.2

*Grain_246:
XU_246 in out fe_tanh Vc=0.44265818498827325 Qo=1.5607732444879095e-13 K=2.62 tau=1.1412158330003126e-07 off=-0.2

*Grain_247:
XU_247 in out fe_tanh Vc=0.7686720607803912 Qo=2.7102690675045385e-13 K=2.62 tau=9.686175526944945e-08 off=-0.2

*Grain_248:
XU_248 in out fe_tanh Vc=0.400667240657868 Qo=1.412716923280579e-13 K=2.62 tau=9.793955638757724e-08 off=-0.2

*Grain_249:
XU_249 in out fe_tanh Vc=-0.21718987407601903 Qo=7.657921076067507e-14 K=2.62 tau=8.995445706272409e-08 off=-0.2

*Grain_250:
XU_250 in out fe_tanh Vc=0.4550267288519956 Qo=1.6043836260202976e-13 K=2.62 tau=8.896357313117196e-08 off=-0.2

*Grain_251:
XU_251 in out fe_tanh Vc=0.5347603360364468 Qo=1.8855172071903764e-13 K=2.62 tau=7.572820312262096e-08 off=-0.2

*Grain_252:
XU_252 in out fe_tanh Vc=0.7283018656196343 Qo=2.5679273631862647e-13 K=2.62 tau=9.756710184583177e-08 off=-0.2

*Grain_253:
XU_253 in out fe_tanh Vc=-0.13170235516811984 Qo=4.6437074734739404e-14 K=2.62 tau=1.1515679470906826e-07 off=-0.2

*Grain_254:
XU_254 in out fe_tanh Vc=0.6569189160189721 Qo=2.3162374551993737e-13 K=2.62 tau=1.1453928276440473e-07 off=-0.2

*Grain_255:
XU_255 in out fe_tanh Vc=0.8215947492148448 Qo=2.896869742553737e-13 K=2.62 tau=9.087363196682147e-08 off=-0.2

*Grain_256:
XU_256 in out fe_tanh Vc=0.6960924925485811 Qo=2.4543599890455127e-13 K=2.62 tau=1.1812991719744538e-07 off=-0.2

*Grain_257:
XU_257 in out fe_tanh Vc=0.4962402593210359 Qo=1.749698855351637e-13 K=2.62 tau=1.0073319277853653e-07 off=-0.2

*Grain_258:
XU_258 in out fe_tanh Vc=0.7457613669739132 Qo=2.6294880063642074e-13 K=2.62 tau=8.720043333840214e-08 off=-0.2

*Grain_259:
XU_259 in out fe_tanh Vc=0.4898718894336492 Qo=1.727244551628553e-13 K=2.62 tau=8.21221768184797e-08 off=-0.2

*Grain_260:
XU_260 in out fe_tanh Vc=0.7383338372533409 Qo=2.6032991996197547e-13 K=2.62 tau=1.0104110658778033e-07 off=-0.2

*Grain_261:
XU_261 in out fe_tanh Vc=0.35049774653715465 Qo=1.2358237656059338e-13 K=2.62 tau=9.893461107567407e-08 off=-0.2

*Grain_262:
XU_262 in out fe_tanh Vc=0.4101904020008906 Qo=1.4462947400502495e-13 K=2.62 tau=9.475690154537733e-08 off=-0.2

*Grain_263:
XU_263 in out fe_tanh Vc=0.570710470707221 Qo=2.0122741727966217e-13 K=2.62 tau=8.356217249089263e-08 off=-0.2

*Grain_264:
XU_264 in out fe_tanh Vc=0.22864992914387464 Qo=8.0619923874506e-14 K=2.62 tau=9.799181030909889e-08 off=-0.2

*Grain_265:
XU_265 in out fe_tanh Vc=0.4948747022966868 Qo=1.7448840231860844e-13 K=2.62 tau=8.612100277795983e-08 off=-0.2

*Grain_266:
XU_266 in out fe_tanh Vc=0.723724441178393 Qo=2.551787773229866e-13 K=2.62 tau=9.883413133438283e-08 off=-0.2

*Grain_267:
XU_267 in out fe_tanh Vc=0.23812549049495801 Qo=8.396092221923704e-14 K=2.62 tau=9.610931616442081e-08 off=-0.2

*Grain_268:
XU_268 in out fe_tanh Vc=0.3593201265905256 Qo=1.266930690106539e-13 K=2.62 tau=8.991276646742397e-08 off=-0.2

*Grain_269:
XU_269 in out fe_tanh Vc=0.5683752641087678 Qo=2.0040404427927048e-13 K=2.62 tau=1.1682535885043592e-07 off=-0.2

*Grain_270:
XU_270 in out fe_tanh Vc=0.5752966502874802 Qo=2.0284446325916326e-13 K=2.62 tau=9.904728568173713e-08 off=-0.2

*Grain_271:
XU_271 in out fe_tanh Vc=0.5933734792011252 Qo=2.0921819176355088e-13 K=2.62 tau=9.282779140140997e-08 off=-0.2

*Grain_272:
XU_272 in out fe_tanh Vc=0.18503859282837842 Qo=6.524295600495365e-14 K=2.62 tau=9.945594234391981e-08 off=-0.2

*Grain_273:
XU_273 in out fe_tanh Vc=-0.05812873939402813 Qo=2.049567459921992e-14 K=2.62 tau=1.0189901902100089e-07 off=-0.2

*Grain_274:
XU_274 in out fe_tanh Vc=0.39253617867104396 Qo=1.384047524569147e-13 K=2.62 tau=8.700923295058768e-08 off=-0.2

*Grain_275:
XU_275 in out fe_tanh Vc=0.7474577150289824 Qo=2.6354691781745994e-13 K=2.62 tau=8.321186800184246e-08 off=-0.2

*Grain_276:
XU_276 in out fe_tanh Vc=0.331566625124619 Qo=1.1690743214730516e-13 K=2.62 tau=9.797516626069846e-08 off=-0.2

*Grain_277:
XU_277 in out fe_tanh Vc=0.19796136929451952 Qo=6.979941162621033e-14 K=2.62 tau=1.010534453306769e-07 off=-0.2

*Grain_278:
XU_278 in out fe_tanh Vc=0.13392629562607178 Qo=4.7221216287255256e-14 K=2.62 tau=1.0151517805346918e-07 off=-0.2

*Grain_279:
XU_279 in out fe_tanh Vc=0.4177774176432644 Qo=1.4730458799177797e-13 K=2.62 tau=1.0399323979331151e-07 off=-0.2

*Grain_280:
XU_280 in out fe_tanh Vc=0.5755575802041595 Qo=2.0293646481848158e-13 K=2.62 tau=1.04293313458143e-07 off=-0.2

*Grain_281:
XU_281 in out fe_tanh Vc=0.6996224758076108 Qo=2.466806394897762e-13 K=2.62 tau=1.0896507125128923e-07 off=-0.2

*Grain_282:
XU_282 in out fe_tanh Vc=0.8356316092027347 Qo=2.9463624578105485e-13 K=2.62 tau=8.428782088907104e-08 off=-0.2

*Grain_283:
XU_283 in out fe_tanh Vc=0.32507479907863346 Qo=1.1461847223555916e-13 K=2.62 tau=1.1267923161935609e-07 off=-0.2

*Grain_284:
XU_284 in out fe_tanh Vc=0.13033001283072349 Qo=4.5953199077375694e-14 K=2.62 tau=1.0286161119989556e-07 off=-0.2

*Grain_285:
XU_285 in out fe_tanh Vc=0.2493579657495214 Qo=8.79213927224899e-14 K=2.62 tau=9.460111933709051e-08 off=-0.2

*Grain_286:
XU_286 in out fe_tanh Vc=0.46989914404241995 Qo=1.6568224343318277e-13 K=2.62 tau=1.0503213265135743e-07 off=-0.2

*Grain_287:
XU_287 in out fe_tanh Vc=0.7134633760299254 Qo=2.515608173514343e-13 K=2.62 tau=9.740312230086465e-08 off=-0.2

*Grain_288:
XU_288 in out fe_tanh Vc=0.7280311152301551 Qo=2.566972721482655e-13 K=2.62 tau=1.0834362729958924e-07 off=-0.2

*Grain_289:
XU_289 in out fe_tanh Vc=0.33757208373039954 Qo=1.1902490324140233e-13 K=2.62 tau=8.921713698348752e-08 off=-0.2

*Grain_290:
XU_290 in out fe_tanh Vc=0.2150642441999452 Qo=7.582973264171789e-14 K=2.62 tau=9.298862189809976e-08 off=-0.2

*Grain_291:
XU_291 in out fe_tanh Vc=0.41906190118230746 Qo=1.4775748542115154e-13 K=2.62 tau=8.797752680313418e-08 off=-0.2

*Grain_292:
XU_292 in out fe_tanh Vc=0.2905433259423435 Qo=1.0244298306770334e-13 K=2.62 tau=1.0378001466527574e-07 off=-0.2

*Grain_293:
XU_293 in out fe_tanh Vc=0.2412672811416681 Qo=8.506868955472579e-14 K=2.62 tau=9.804251887588834e-08 off=-0.2

*Grain_294:
XU_294 in out fe_tanh Vc=0.3923948218337669 Qo=1.383549112979732e-13 K=2.62 tau=1.0413487283481522e-07 off=-0.2

*Grain_295:
XU_295 in out fe_tanh Vc=0.7584333119358428 Qo=2.6741681530844743e-13 K=2.62 tau=9.867279452120401e-08 off=-0.2

*Grain_296:
XU_296 in out fe_tanh Vc=0.5319546098447834 Qo=1.8756244671037489e-13 K=2.62 tau=1.1082086578435771e-07 off=-0.2

*Grain_297:
XU_297 in out fe_tanh Vc=0.22898777277690993 Qo=8.073904452360822e-14 K=2.62 tau=8.915432569081254e-08 off=-0.2

*Grain_298:
XU_298 in out fe_tanh Vc=0.7350245415102561 Qo=2.591630918248111e-13 K=2.62 tau=9.821058950005949e-08 off=-0.2

*Grain_299:
XU_299 in out fe_tanh Vc=0.7242964629114095 Qo=2.5538046707965096e-13 K=2.62 tau=9.871144029716946e-08 off=-0.2

*Grain_300:
XU_300 in out fe_tanh Vc=0.4359483856422091 Qo=1.5371150909726939e-13 K=2.62 tau=1.024250955823657e-07 off=-0.2

*Grain_301:
XU_301 in out fe_tanh Vc=0.6259660331832031 Qo=2.2071003534622467e-13 K=2.62 tau=1.0294750460044324e-07 off=-0.2

*Grain_302:
XU_302 in out fe_tanh Vc=0.3770489040664202 Qo=1.3294407768512116e-13 K=2.62 tau=8.627419419663537e-08 off=-0.2

*Grain_303:
XU_303 in out fe_tanh Vc=0.18896174697178386 Qo=6.662622513420094e-14 K=2.62 tau=1.1645881179838197e-07 off=-0.2

*Grain_304:
XU_304 in out fe_tanh Vc=0.5065809596034238 Qo=1.7861592414403909e-13 K=2.62 tau=1.0791065524035906e-07 off=-0.2

*Grain_305:
XU_305 in out fe_tanh Vc=0.2039639598506845 Qo=7.191587147161596e-14 K=2.62 tau=8.997410077370851e-08 off=-0.2

*Grain_306:
XU_306 in out fe_tanh Vc=0.41218256192204306 Qo=1.4533189180935366e-13 K=2.62 tau=1.0759480949013731e-07 off=-0.2

*Grain_307:
XU_307 in out fe_tanh Vc=0.21048628352320542 Qo=7.421558457422817e-14 K=2.62 tau=9.673507809981235e-08 off=-0.2

*Grain_308:
XU_308 in out fe_tanh Vc=-0.2844387864846107 Qo=1.002905769496955e-13 K=2.62 tau=1.1264148687975323e-07 off=-0.2

*Grain_309:
XU_309 in out fe_tanh Vc=0.15987104379502237 Qo=5.636910288470912e-14 K=2.62 tau=1.1201442165573353e-07 off=-0.2

*Grain_310:
XU_310 in out fe_tanh Vc=0.3369745058291024 Qo=1.188142026079403e-13 K=2.62 tau=9.270769745575022e-08 off=-0.2

*Grain_311:
XU_311 in out fe_tanh Vc=0.4458353474761531 Qo=1.5719756357971426e-13 K=2.62 tau=1.0309108350075091e-07 off=-0.2

*Grain_312:
XU_312 in out fe_tanh Vc=0.6297363018399196 Qo=2.2203939841766328e-13 K=2.62 tau=1.1154067845303822e-07 off=-0.2

*Grain_313:
XU_313 in out fe_tanh Vc=0.21179437230170203 Qo=7.467680500031078e-14 K=2.62 tau=1.1406039619375716e-07 off=-0.2

*Grain_314:
XU_314 in out fe_tanh Vc=0.8161706873844472 Qo=2.87774498474189e-13 K=2.62 tau=9.926552192775101e-08 off=-0.2

*Grain_315:
XU_315 in out fe_tanh Vc=0.1945778242549765 Qo=6.860640384993293e-14 K=2.62 tau=1.173955206644147e-07 off=-0.2

*Grain_316:
XU_316 in out fe_tanh Vc=0.5673189163442619 Qo=2.0003158548744692e-13 K=2.62 tau=1.1481318505931197e-07 off=-0.2

*Grain_317:
XU_317 in out fe_tanh Vc=0.06504223926556102 Qo=2.293331293760171e-14 K=2.62 tau=9.812734058512688e-08 off=-0.2

*Grain_318:
XU_318 in out fe_tanh Vc=0.2993581855473991 Qo=1.055510238748224e-13 K=2.62 tau=1.1014855176487026e-07 off=-0.2

*Grain_319:
XU_319 in out fe_tanh Vc=0.7229757197099862 Qo=2.549147848170095e-13 K=2.62 tau=1.0592305913121581e-07 off=-0.2

*Grain_320:
XU_320 in out fe_tanh Vc=0.8168180257257167 Qo=2.8800274419457737e-13 K=2.62 tau=1.0473732003742723e-07 off=-0.2

*Grain_321:
XU_321 in out fe_tanh Vc=0.6997710757453964 Qo=2.467330345012983e-13 K=2.62 tau=9.586151661389292e-08 off=-0.2

*Grain_322:
XU_322 in out fe_tanh Vc=0.2807409047462801 Qo=9.89867368594869e-14 K=2.62 tau=1.0605666842443398e-07 off=-0.2

*Grain_323:
XU_323 in out fe_tanh Vc=0.8726982265758392 Qo=3.0770560417575954e-13 K=2.62 tau=8.922099145900935e-08 off=-0.2

*Grain_324:
XU_324 in out fe_tanh Vc=-0.00821442940367162 Qo=2.896334478108675e-15 K=2.62 tau=1.0256938581151252e-07 off=-0.2

*Grain_325:
XU_325 in out fe_tanh Vc=0.841306729534975 Qo=2.9663724254880795e-13 K=2.62 tau=1.0447020076773996e-07 off=-0.2

*Grain_326:
XU_326 in out fe_tanh Vc=0.12040316163724257 Qo=4.245307996284756e-14 K=2.62 tau=1.0127561864896839e-07 off=-0.2

*Grain_327:
XU_327 in out fe_tanh Vc=0.06971757285994412 Qo=2.4581793826611352e-14 K=2.62 tau=8.848413966871998e-08 off=-0.2

*Grain_328:
XU_328 in out fe_tanh Vc=0.9220808717477404 Qo=3.251174840280174e-13 K=2.62 tau=1.0455467440117582e-07 off=-0.2

*Grain_329:
XU_329 in out fe_tanh Vc=0.2751024860361815 Qo=9.699868075606817e-14 K=2.62 tau=9.494689829308834e-08 off=-0.2

*Grain_330:
XU_330 in out fe_tanh Vc=0.20104458919205948 Qo=7.088652743839861e-14 K=2.62 tau=9.779408025511967e-08 off=-0.2

*Grain_331:
XU_331 in out fe_tanh Vc=0.2534276490143934 Qo=8.935632671191128e-14 K=2.62 tau=1.2911763052693344e-07 off=-0.2

*Grain_332:
XU_332 in out fe_tanh Vc=0.24613827970685667 Qo=8.678616016575419e-14 K=2.62 tau=1.2023193370999147e-07 off=-0.2

*Grain_333:
XU_333 in out fe_tanh Vc=0.4045281934307254 Qo=1.4263302980931714e-13 K=2.62 tau=1.0057253966443989e-07 off=-0.2

*Grain_334:
XU_334 in out fe_tanh Vc=0.22689256720592765 Qo=8.000029374303069e-14 K=2.62 tau=9.901251822521893e-08 off=-0.2

*Grain_335:
XU_335 in out fe_tanh Vc=0.132804386125065 Qo=4.6825641012406444e-14 K=2.62 tau=1.0069643711241403e-07 off=-0.2

*Grain_336:
XU_336 in out fe_tanh Vc=0.3010275060052709 Qo=1.0613961136636321e-13 K=2.62 tau=1.0181616209507467e-07 off=-0.2

*Grain_337:
XU_337 in out fe_tanh Vc=0.30238323605064565 Qo=1.0661762967785684e-13 K=2.62 tau=1.046480436987181e-07 off=-0.2

*Grain_338:
XU_338 in out fe_tanh Vc=0.6252662370150414 Qo=2.2046329346436135e-13 K=2.62 tau=1.0708587124911063e-07 off=-0.2

*Grain_339:
XU_339 in out fe_tanh Vc=0.45502423984557927 Qo=1.6043748500058655e-13 K=2.62 tau=9.75700617709437e-08 off=-0.2

*Grain_340:
XU_340 in out fe_tanh Vc=0.43770026104277454 Qo=1.543292047246419e-13 K=2.62 tau=9.638626374349934e-08 off=-0.2

*Grain_341:
XU_341 in out fe_tanh Vc=0.6559091914458665 Qo=2.3126772564919964e-13 K=2.62 tau=1.0892669438675988e-07 off=-0.2

*Grain_342:
XU_342 in out fe_tanh Vc=0.45779614063141383 Qo=1.6141483247311101e-13 K=2.62 tau=9.287726058456959e-08 off=-0.2

*Grain_343:
XU_343 in out fe_tanh Vc=0.5013458071294619 Qo=1.7677005611555323e-13 K=2.62 tau=1.0320522410116548e-07 off=-0.2

*Grain_344:
XU_344 in out fe_tanh Vc=0.3086409025516814 Qo=1.0882402702437911e-13 K=2.62 tau=1.0095915873658086e-07 off=-0.2

*Grain_345:
XU_345 in out fe_tanh Vc=0.3887197440442917 Qo=1.3705911167656179e-13 K=2.62 tau=8.734933384898697e-08 off=-0.2

*Grain_346:
XU_346 in out fe_tanh Vc=0.20081938482778983 Qo=7.080712238994044e-14 K=2.62 tau=8.76210155730703e-08 off=-0.2

*Grain_347:
XU_347 in out fe_tanh Vc=0.5233175780885337 Qo=1.845171064152883e-13 K=2.62 tau=1.0753854120023986e-07 off=-0.2

*Grain_348:
XU_348 in out fe_tanh Vc=1.1030715750723743 Qo=3.8893319032917187e-13 K=2.62 tau=9.014752268639145e-08 off=-0.2

*Grain_349:
XU_349 in out fe_tanh Vc=0.3148536772598921 Qo=1.1101459592549709e-13 K=2.62 tau=9.896839912175382e-08 off=-0.2

*Grain_350:
XU_350 in out fe_tanh Vc=0.5132069061798289 Qo=1.8095217375752663e-13 K=2.62 tau=8.509369234653561e-08 off=-0.2

*Grain_351:
XU_351 in out fe_tanh Vc=0.4012215817291507 Qo=1.414671480412289e-13 K=2.62 tau=7.403015344507635e-08 off=-0.2

*Grain_352:
XU_352 in out fe_tanh Vc=0.6727814805773227 Qo=2.3721674417922834e-13 K=2.62 tau=9.298559506061162e-08 off=-0.2

*Grain_353:
XU_353 in out fe_tanh Vc=0.669889643076084 Qo=2.361971080915189e-13 K=2.62 tau=1.1761986652782663e-07 off=-0.2

*Grain_354:
XU_354 in out fe_tanh Vc=0.18881719123249635 Qo=6.657525607096694e-14 K=2.62 tau=1.0437286811790565e-07 off=-0.2

*Grain_355:
XU_355 in out fe_tanh Vc=0.6839286192142038 Qo=2.4114712575288036e-13 K=2.62 tau=9.481545255921712e-08 off=-0.2

*Grain_356:
XU_356 in out fe_tanh Vc=0.32589462452443885 Qo=1.149075353692268e-13 K=2.62 tau=9.401370643124966e-08 off=-0.2

*Grain_357:
XU_357 in out fe_tanh Vc=0.7165691780178957 Qo=2.5265589540711955e-13 K=2.62 tau=1.1497809034518841e-07 off=-0.2

*Grain_358:
XU_358 in out fe_tanh Vc=0.8607644926037584 Qo=3.0349787610879664e-13 K=2.62 tau=1.0250958980883679e-07 off=-0.2

*Grain_359:
XU_359 in out fe_tanh Vc=0.09706475549805349 Qo=3.4224166298458025e-14 K=2.62 tau=1.1161752008417674e-07 off=-0.2

*Grain_360:
XU_360 in out fe_tanh Vc=0.7062152018597223 Qo=2.49005175842955e-13 K=2.62 tau=1.008918381665144e-07 off=-0.2

*Grain_361:
XU_361 in out fe_tanh Vc=0.5360337816195886 Qo=1.8900072626369544e-13 K=2.62 tau=9.452660546456175e-08 off=-0.2

*Grain_362:
XU_362 in out fe_tanh Vc=0.2788033454893649 Qo=9.830357076195202e-14 K=2.62 tau=1.0910636949182382e-07 off=-0.2

*Grain_363:
XU_363 in out fe_tanh Vc=0.07760095569401781 Qo=2.7361404239508937e-14 K=2.62 tau=1.184355812850462e-07 off=-0.2

*Grain_364:
XU_364 in out fe_tanh Vc=0.1621832836214505 Qo=5.718437800630751e-14 K=2.62 tau=1.0321462945395966e-07 off=-0.2

*Grain_365:
XU_365 in out fe_tanh Vc=-0.0888636784714329 Qo=3.133253974930183e-14 K=2.62 tau=9.381687826012269e-08 off=-0.2

*Grain_366:
XU_366 in out fe_tanh Vc=1.2634156181290759 Qo=4.4546906853111837e-13 K=2.62 tau=1.0534382342023566e-07 off=-0.2

*Grain_367:
XU_367 in out fe_tanh Vc=0.6920417713931144 Qo=2.4400775078563286e-13 K=2.62 tau=8.40468243167349e-08 off=-0.2

*Grain_368:
XU_368 in out fe_tanh Vc=0.752887739572899 Qo=2.6546149599820276e-13 K=2.62 tau=1.1957331303887818e-07 off=-0.2

*Grain_369:
XU_369 in out fe_tanh Vc=-0.17041778024681992 Qo=6.008778800764817e-14 K=2.62 tau=1.0740720451500833e-07 off=-0.2

*Grain_370:
XU_370 in out fe_tanh Vc=0.4740868636776314 Qo=1.6715879599308358e-13 K=2.62 tau=9.515511969168126e-08 off=-0.2

*Grain_371:
XU_371 in out fe_tanh Vc=0.27664927470222933 Qo=9.754406463164443e-14 K=2.62 tau=1.0881450923338383e-07 off=-0.2

*Grain_372:
XU_372 in out fe_tanh Vc=0.4517615709783748 Qo=1.5928709708362275e-13 K=2.62 tau=1.1915594155265067e-07 off=-0.2

*Grain_373:
XU_373 in out fe_tanh Vc=1.0770222107322291 Qo=3.797484170036559e-13 K=2.62 tau=1.1005430752177602e-07 off=-0.2

*Grain_374:
XU_374 in out fe_tanh Vc=0.6592222781585154 Qo=2.324358904483907e-13 K=2.62 tau=1.0481578477281293e-07 off=-0.2

*Grain_375:
XU_375 in out fe_tanh Vc=0.49801214964322565 Qo=1.7559463824522916e-13 K=2.62 tau=1.2729518032274393e-07 off=-0.2

*Grain_376:
XU_376 in out fe_tanh Vc=0.4610505417316571 Qo=1.6256230524925006e-13 K=2.62 tau=1.0746233903941177e-07 off=-0.2

*Grain_377:
XU_377 in out fe_tanh Vc=0.6573386538144034 Qo=2.3177174131963706e-13 K=2.62 tau=1.0790645750536487e-07 off=-0.2

*Grain_378:
XU_378 in out fe_tanh Vc=0.8017087561278584 Qo=2.8267535061374555e-13 K=2.62 tau=9.307813889305726e-08 off=-0.2

*Grain_379:
XU_379 in out fe_tanh Vc=0.3490281131399507 Qo=1.2306419694405187e-13 K=2.62 tau=1.0110343288066077e-07 off=-0.2

*Grain_380:
XU_380 in out fe_tanh Vc=0.3537011880735629 Qo=1.247118814494366e-13 K=2.62 tau=1.0162226925522461e-07 off=-0.2

*Grain_381:
XU_381 in out fe_tanh Vc=0.289991056188461 Qo=1.0224825768255711e-13 K=2.62 tau=1.168309950098073e-07 off=-0.2

*Grain_382:
XU_382 in out fe_tanh Vc=0.08043958509361804 Qo=2.83622796255656e-14 K=2.62 tau=9.372784344461182e-08 off=-0.2

*Grain_383:
XU_383 in out fe_tanh Vc=0.5073920301664887 Qo=1.7890190038420668e-13 K=2.62 tau=1.0748010527337466e-07 off=-0.2

*Grain_384:
XU_384 in out fe_tanh Vc=0.3801968851977124 Qo=1.3405402773021152e-13 K=2.62 tau=1.0694979270505085e-07 off=-0.2

*Grain_385:
XU_385 in out fe_tanh Vc=0.07205665577911469 Qo=2.5406533583084356e-14 K=2.62 tau=1.1474891377016883e-07 off=-0.2

*Grain_386:
XU_386 in out fe_tanh Vc=0.3131838660181739 Qo=1.1042583538795321e-13 K=2.62 tau=1.1588616112211539e-07 off=-0.2

*Grain_387:
XU_387 in out fe_tanh Vc=0.2852800234551003 Qo=1.0058718959582764e-13 K=2.62 tau=1.1418429889370222e-07 off=-0.2

*Grain_388:
XU_388 in out fe_tanh Vc=0.3668879094741414 Qo=1.293614016983583e-13 K=2.62 tau=1.1250448099439624e-07 off=-0.2

*Grain_389:
XU_389 in out fe_tanh Vc=-0.09659908099804343 Qo=3.4059973626797555e-14 K=2.62 tau=8.564952127175051e-08 off=-0.2

*Grain_390:
XU_390 in out fe_tanh Vc=0.9711485392635546 Qo=3.42418305570522e-13 K=2.62 tau=8.477742235432443e-08 off=-0.2

*Grain_391:
XU_391 in out fe_tanh Vc=0.7347453026768143 Qo=2.590646347048846e-13 K=2.62 tau=7.517713579829263e-08 off=-0.2

*Grain_392:
XU_392 in out fe_tanh Vc=0.9584472655214091 Qo=3.379399498324072e-13 K=2.62 tau=9.578503691050523e-08 off=-0.2

*Grain_393:
XU_393 in out fe_tanh Vc=0.6464453758811546 Qo=2.279308687638894e-13 K=2.62 tau=7.902181707355828e-08 off=-0.2

*Grain_394:
XU_394 in out fe_tanh Vc=0.5070239049966758 Qo=1.787721027355578e-13 K=2.62 tau=1.095184593932857e-07 off=-0.2

*Grain_395:
XU_395 in out fe_tanh Vc=0.22368533203718785 Qo=7.886945125329285e-14 K=2.62 tau=9.294503378217019e-08 off=-0.2

*Grain_396:
XU_396 in out fe_tanh Vc=0.40188322964008205 Qo=1.4170043918813958e-13 K=2.62 tau=9.0517907745579e-08 off=-0.2

*Grain_397:
XU_397 in out fe_tanh Vc=0.44432254874024674 Qo=1.566641642500802e-13 K=2.62 tau=1.0511894444017032e-07 off=-0.2

*Grain_398:
XU_398 in out fe_tanh Vc=0.8879016971286018 Qo=3.1306621217236537e-13 K=2.62 tau=1.0464086932008556e-07 off=-0.2

*Grain_399:
XU_399 in out fe_tanh Vc=-0.062124737168809674 Qo=2.1904627742620508e-14 K=2.62 tau=9.239761313197357e-08 off=-0.2

*Grain_400:
XU_400 in out fe_tanh Vc=0.3195324885168319 Qo=1.1266430300727939e-13 K=2.62 tau=8.646433974692629e-08 off=-0.2

*Grain_401:
XU_401 in out fe_tanh Vc=0.7725195615430508 Qo=2.723835011730025e-13 K=2.62 tau=8.678554499785248e-08 off=-0.2

*Grain_402:
XU_402 in out fe_tanh Vc=0.462935746689417 Qo=1.632270116882659e-13 K=2.62 tau=1.038204050276372e-07 off=-0.2

*Grain_403:
XU_403 in out fe_tanh Vc=0.3135034418021565 Qo=1.1053851495655524e-13 K=2.62 tau=9.788502771732814e-08 off=-0.2

*Grain_404:
XU_404 in out fe_tanh Vc=0.41646414883772587 Qo=1.468415411344021e-13 K=2.62 tau=9.352435306321164e-08 off=-0.2

*Grain_405:
XU_405 in out fe_tanh Vc=0.4293118919502608 Qo=1.513715406649947e-13 K=2.62 tau=8.494903855412874e-08 off=-0.2

*Grain_406:
XU_406 in out fe_tanh Vc=0.8812222622698438 Qo=3.107111030680063e-13 K=2.62 tau=8.476587790969025e-08 off=-0.2

*Grain_407:
XU_407 in out fe_tanh Vc=0.586875138618104 Qo=2.0692693488420096e-13 K=2.62 tau=9.993842734602585e-08 off=-0.2

*Grain_408:
XU_408 in out fe_tanh Vc=0.5569321642518749 Qo=1.9636930942146702e-13 K=2.62 tau=8.711931475588843e-08 off=-0.2

*Grain_409:
XU_409 in out fe_tanh Vc=-0.16916027674325546 Qo=5.964440349793551e-14 K=2.62 tau=1.0506323761503604e-07 off=-0.2

*Grain_410:
XU_410 in out fe_tanh Vc=0.2948929975348483 Qo=1.039766384420122e-13 K=2.62 tau=8.097547847290589e-08 off=-0.2

*Grain_411:
XU_411 in out fe_tanh Vc=0.6553530946481072 Qo=2.3107165088254627e-13 K=2.62 tau=9.123170563935521e-08 off=-0.2

*Grain_412:
XU_412 in out fe_tanh Vc=0.09145903430388413 Qo=3.224763904726756e-14 K=2.62 tau=8.338002700114084e-08 off=-0.2

*Grain_413:
XU_413 in out fe_tanh Vc=0.582641822814004 Qo=2.054343055221838e-13 K=2.62 tau=1.013131246964434e-07 off=-0.2

*Grain_414:
XU_414 in out fe_tanh Vc=0.804913601327881 Qo=2.838053504218488e-13 K=2.62 tau=9.378755534167105e-08 off=-0.2

*Grain_415:
XU_415 in out fe_tanh Vc=0.5866234613200152 Qo=2.0683819571560012e-13 K=2.62 tau=9.14313489058395e-08 off=-0.2

*Grain_416:
XU_416 in out fe_tanh Vc=0.5332948198528895 Qo=1.8803499279527384e-13 K=2.62 tau=9.839358927113928e-08 off=-0.2

*Grain_417:
XU_417 in out fe_tanh Vc=0.35926188559976097 Qo=1.2667253375722346e-13 K=2.62 tau=1.0541315211042676e-07 off=-0.2

*Grain_418:
XU_418 in out fe_tanh Vc=0.5985518193481563 Qo=2.1104402827272056e-13 K=2.62 tau=9.33247095542275e-08 off=-0.2

*Grain_419:
XU_419 in out fe_tanh Vc=0.3163726673351128 Qo=1.1155017826610377e-13 K=2.62 tau=9.163242242748658e-08 off=-0.2

*Grain_420:
XU_420 in out fe_tanh Vc=0.5838532617147227 Qo=2.0586144806414846e-13 K=2.62 tau=8.134994020333488e-08 off=-0.2

*Grain_421:
XU_421 in out fe_tanh Vc=0.07566851920116707 Qo=2.6680044382852636e-14 K=2.62 tau=1.0428590593309646e-07 off=-0.2

*Grain_422:
XU_422 in out fe_tanh Vc=0.579547531289842 Qo=2.0434328595328423e-13 K=2.62 tau=8.545517145234644e-08 off=-0.2

*Grain_423:
XU_423 in out fe_tanh Vc=0.7560090867370652 Qo=2.6656205514424405e-13 K=2.62 tau=9.676593105850663e-08 off=-0.2

*Grain_424:
XU_424 in out fe_tanh Vc=0.06335990566029082 Qo=2.2340137126455653e-14 K=2.62 tau=8.188341689589778e-08 off=-0.2

*Grain_425:
XU_425 in out fe_tanh Vc=0.8680102113612977 Qo=3.0605265186069e-13 K=2.62 tau=9.448342845380643e-08 off=-0.2

*Grain_426:
XU_426 in out fe_tanh Vc=0.9705544453177484 Qo=3.4220883334866505e-13 K=2.62 tau=1.2003533526047513e-07 off=-0.2

*Grain_427:
XU_427 in out fe_tanh Vc=0.4593452336571035 Qo=1.6196102884532615e-13 K=2.62 tau=9.322393811361086e-08 off=-0.2

*Grain_428:
XU_428 in out fe_tanh Vc=0.13376664765744817 Qo=4.716492583868461e-14 K=2.62 tau=9.663693672443922e-08 off=-0.2

*Grain_429:
XU_429 in out fe_tanh Vc=0.4037226290713393 Qo=1.4234899500741323e-13 K=2.62 tau=9.513096828251198e-08 off=-0.2

*Grain_430:
XU_430 in out fe_tanh Vc=0.4207856355593479 Qo=1.48365258774842e-13 K=2.62 tau=9.833963571799572e-08 off=-0.2

*Grain_431:
XU_431 in out fe_tanh Vc=0.6117967520166679 Qo=2.1571407329506764e-13 K=2.62 tau=1.0062504391751816e-07 off=-0.2

*Grain_432:
XU_432 in out fe_tanh Vc=0.5517297802460914 Qo=1.9453499526233908e-13 K=2.62 tau=9.846780539958845e-08 off=-0.2

*Grain_433:
XU_433 in out fe_tanh Vc=0.9063717286958304 Qo=3.195785804223145e-13 K=2.62 tau=1.1638905235961424e-07 off=-0.2

*Grain_434:
XU_434 in out fe_tanh Vc=0.42773480276906145 Qo=1.5081547309826656e-13 K=2.62 tau=1.0811004012739085e-07 off=-0.2

*Grain_435:
XU_435 in out fe_tanh Vc=0.7449777300519103 Qo=2.6267249725319346e-13 K=2.62 tau=1.0004342461083075e-07 off=-0.2

*Grain_436:
XU_436 in out fe_tanh Vc=0.0745301463170196 Qo=2.627866426607585e-14 K=2.62 tau=1.0540455132295566e-07 off=-0.2

*Grain_437:
XU_437 in out fe_tanh Vc=0.12430138770386873 Qo=4.3827559674753626e-14 K=2.62 tau=9.353535012049701e-08 off=-0.2

*Grain_438:
XU_438 in out fe_tanh Vc=0.3890658839384005 Qo=1.371811575132584e-13 K=2.62 tau=9.622840308840181e-08 off=-0.2

*Grain_439:
XU_439 in out fe_tanh Vc=0.282262499826966 Qo=9.952323770176588e-14 K=2.62 tau=1.0380987168622531e-07 off=-0.2

*Grain_440:
XU_440 in out fe_tanh Vc=0.5198205178358916 Qo=1.8328407418821432e-13 K=2.62 tau=1.1215397583018337e-07 off=-0.2

*Grain_441:
XU_441 in out fe_tanh Vc=0.6212303180835972 Qo=2.1904026447749485e-13 K=2.62 tau=8.890136578077613e-08 off=-0.2

*Grain_442:
XU_442 in out fe_tanh Vc=0.13672870538500193 Qo=4.82093209513418e-14 K=2.62 tau=9.485376403909497e-08 off=-0.2

*Grain_443:
XU_443 in out fe_tanh Vc=0.5565813850872724 Qo=1.962456278194088e-13 K=2.62 tau=9.037532713846812e-08 off=-0.2

*Grain_444:
XU_444 in out fe_tanh Vc=0.3317311137016319 Qo=1.1696542935118208e-13 K=2.62 tau=1.1475474041134549e-07 off=-0.2

*Grain_445:
XU_445 in out fe_tanh Vc=0.5719699921046896 Qo=2.0167151328075182e-13 K=2.62 tau=9.803916313275994e-08 off=-0.2

*Grain_446:
XU_446 in out fe_tanh Vc=0.9249965098096466 Qo=3.261455119809523e-13 K=2.62 tau=1.1244941441694208e-07 off=-0.2

*Grain_447:
XU_447 in out fe_tanh Vc=0.3171969276901551 Qo=1.1184080510917822e-13 K=2.62 tau=1.1175232505806663e-07 off=-0.2

*Grain_448:
XU_448 in out fe_tanh Vc=0.4227932855361554 Qo=1.4907313823451607e-13 K=2.62 tau=8.496262951472307e-08 off=-0.2

*Grain_449:
XU_449 in out fe_tanh Vc=0.45994113220948146 Qo=1.621711373553507e-13 K=2.62 tau=9.259508479044762e-08 off=-0.2

*Grain_450:
XU_450 in out fe_tanh Vc=-0.5782732293155302 Qo=2.0389397845274477e-13 K=2.62 tau=1.2659084928724185e-07 off=-0.2

*Grain_451:
XU_451 in out fe_tanh Vc=0.30632324105264835 Qo=1.080068402694191e-13 K=2.62 tau=1.0223669608817688e-07 off=-0.2

*Grain_452:
XU_452 in out fe_tanh Vc=0.45361872524762165 Qo=1.5994191310027533e-13 K=2.62 tau=9.871089953199174e-08 off=-0.2

*Grain_453:
XU_453 in out fe_tanh Vc=-0.05577178857934023 Qo=1.9664634782292938e-14 K=2.62 tau=1.001552566439474e-07 off=-0.2

*Grain_454:
XU_454 in out fe_tanh Vc=0.7261602946923653 Qo=2.5603763752732244e-13 K=2.62 tau=9.751653632116404e-08 off=-0.2

*Grain_455:
XU_455 in out fe_tanh Vc=0.7279640449240665 Qo=2.566736237570705e-13 K=2.62 tau=9.879970635563502e-08 off=-0.2

*Grain_456:
XU_456 in out fe_tanh Vc=0.34727867863627 Qo=1.2244736195513121e-13 K=2.62 tau=1.1077417737300383e-07 off=-0.2

*Grain_457:
XU_457 in out fe_tanh Vc=0.31816827050787616 Qo=1.1218329191559853e-13 K=2.62 tau=9.694708418661985e-08 off=-0.2

*Grain_458:
XU_458 in out fe_tanh Vc=0.4605679581521704 Qo=1.6239215058711227e-13 K=2.62 tau=1.2348732984340373e-07 off=-0.2

*Grain_459:
XU_459 in out fe_tanh Vc=0.4818150057077388 Qo=1.698836698843262e-13 K=2.62 tau=9.851400940550618e-08 off=-0.2

*Grain_460:
XU_460 in out fe_tanh Vc=0.8058889221010326 Qo=2.8414923981984304e-13 K=2.62 tau=1.0918054619337243e-07 off=-0.2

*Grain_461:
XU_461 in out fe_tanh Vc=0.3726653054945952 Qo=1.3139845996076774e-13 K=2.62 tau=9.777247167476452e-08 off=-0.2

*Grain_462:
XU_462 in out fe_tanh Vc=0.26926374365291506 Qo=9.493999231376562e-14 K=2.62 tau=1.119300065362711e-07 off=-0.2

*Grain_463:
XU_463 in out fe_tanh Vc=0.3324908655423663 Qo=1.172333110679745e-13 K=2.62 tau=1.0474048455489391e-07 off=-0.2

*Grain_464:
XU_464 in out fe_tanh Vc=0.4331647327447676 Qo=1.5273001793510258e-13 K=2.62 tau=9.786271524845514e-08 off=-0.2

*Grain_465:
XU_465 in out fe_tanh Vc=1.068591892259363 Qo=3.767759619669755e-13 K=2.62 tau=8.333103262560877e-08 off=-0.2

*Grain_466:
XU_466 in out fe_tanh Vc=0.6072873951071345 Qo=2.1412411430347394e-13 K=2.62 tau=1.1700100671504758e-07 off=-0.2

*Grain_467:
XU_467 in out fe_tanh Vc=0.5277473563713596 Qo=1.860790066934976e-13 K=2.62 tau=1.0480686548274775e-07 off=-0.2

*Grain_468:
XU_468 in out fe_tanh Vc=0.6933663408329465 Qo=2.444747821457806e-13 K=2.62 tau=8.337141640972336e-08 off=-0.2

*Grain_469:
XU_469 in out fe_tanh Vc=0.14631373760164523 Qo=5.158891774603065e-14 K=2.62 tau=1.0188347738415837e-07 off=-0.2

*Grain_470:
XU_470 in out fe_tanh Vc=0.4794492345856545 Qo=1.6904952010574953e-13 K=2.62 tau=1.1101266453179046e-07 off=-0.2

*Grain_471:
XU_471 in out fe_tanh Vc=0.5525912799386135 Qo=1.9483875236337597e-13 K=2.62 tau=1.1421611679141924e-07 off=-0.2

*Grain_472:
XU_472 in out fe_tanh Vc=0.2735468439155433 Qo=9.645017523143751e-14 K=2.62 tau=8.688456463561959e-08 off=-0.2

*Grain_473:
XU_473 in out fe_tanh Vc=0.2878181558689946 Qo=1.0148211242723958e-13 K=2.62 tau=1.2451738516179322e-07 off=-0.2

*Grain_474:
XU_474 in out fe_tanh Vc=0.32293996796598945 Qo=1.138657498427261e-13 K=2.62 tau=1.144896257216139e-07 off=-0.2

*Grain_475:
XU_475 in out fe_tanh Vc=0.5270863759749488 Qo=1.8584595090624805e-13 K=2.62 tau=9.177156972342812e-08 off=-0.2

*Grain_476:
XU_476 in out fe_tanh Vc=0.3042364927358203 Qo=1.0727107144115907e-13 K=2.62 tau=9.97084472598575e-08 off=-0.2

*Grain_477:
XU_477 in out fe_tanh Vc=0.07848132797631624 Qo=2.767181564722673e-14 K=2.62 tau=1.0357218431781931e-07 off=-0.2

*Grain_478:
XU_478 in out fe_tanh Vc=-0.020958529815149785 Qo=7.38979051751963e-15 K=2.62 tau=1.0367540051330872e-07 off=-0.2

*Grain_479:
XU_479 in out fe_tanh Vc=0.6274904639924891 Qo=2.2124753604109368e-13 K=2.62 tau=9.967161832338627e-08 off=-0.2

*Grain_480:
XU_480 in out fe_tanh Vc=0.926377748284658 Qo=3.2663252433702386e-13 K=2.62 tau=1.0441471841977256e-07 off=-0.2

*Grain_481:
XU_481 in out fe_tanh Vc=0.3812174930095326 Qo=1.3441388493376616e-13 K=2.62 tau=9.639785932786343e-08 off=-0.2

*Grain_482:
XU_482 in out fe_tanh Vc=0.22605732909447165 Qo=7.97057962410424e-14 K=2.62 tau=9.16183813361762e-08 off=-0.2

*Grain_483:
XU_483 in out fe_tanh Vc=0.6055382552858599 Qo=2.1350738321693909e-13 K=2.62 tau=1.0582924518073333e-07 off=-0.2

*Grain_484:
XU_484 in out fe_tanh Vc=0.8854974233521551 Qo=3.1221848670157097e-13 K=2.62 tau=9.969444091493229e-08 off=-0.2

*Grain_485:
XU_485 in out fe_tanh Vc=0.2688043965934438 Qo=9.477803064115453e-14 K=2.62 tau=1.1456428782901845e-07 off=-0.2

*Grain_486:
XU_486 in out fe_tanh Vc=0.6210154625161535 Qo=2.1896450832241452e-13 K=2.62 tau=1.0508334790742685e-07 off=-0.2

*Grain_487:
XU_487 in out fe_tanh Vc=0.000924169665680652 Qo=3.258539741222474e-16 K=2.62 tau=1.1602077770351244e-07 off=-0.2

*Grain_488:
XU_488 in out fe_tanh Vc=0.2992882766169985 Qo=1.0552637461003519e-13 K=2.62 tau=1.0398840158622563e-07 off=-0.2

*Grain_489:
XU_489 in out fe_tanh Vc=-0.18423549457511984 Qo=6.495979073005555e-14 K=2.62 tau=1.0840154869927829e-07 off=-0.2

*Grain_490:
XU_490 in out fe_tanh Vc=0.4841943979325268 Qo=1.7072262234212163e-13 K=2.62 tau=1.0106361459804344e-07 off=-0.2

*Grain_491:
XU_491 in out fe_tanh Vc=0.46392610549722374 Qo=1.6357620336303606e-13 K=2.62 tau=9.775997031251878e-08 off=-0.2

*Grain_492:
XU_492 in out fe_tanh Vc=0.7236930243210449 Qo=2.551677000195417e-13 K=2.62 tau=1.011416619948551e-07 off=-0.2

*Grain_493:
XU_493 in out fe_tanh Vc=0.3319647266832285 Qo=1.170477992030466e-13 K=2.62 tau=1.046376278519792e-07 off=-0.2

*Grain_494:
XU_494 in out fe_tanh Vc=0.22162711431498233 Qo=7.814374205800613e-14 K=2.62 tau=9.162220453483731e-08 off=-0.2

*Grain_495:
XU_495 in out fe_tanh Vc=0.20564711844131453 Qo=7.25093381652353e-14 K=2.62 tau=9.592095968111715e-08 off=-0.2

*Grain_496:
XU_496 in out fe_tanh Vc=1.0667160047630084 Qo=3.76114540781675e-13 K=2.62 tau=9.998047047612074e-08 off=-0.2

*Grain_497:
XU_497 in out fe_tanh Vc=0.8073135098073888 Qo=2.8465153672791124e-13 K=2.62 tau=1.1509608766326103e-07 off=-0.2

*Grain_498:
XU_498 in out fe_tanh Vc=0.48057998700610416 Qo=1.694482133150538e-13 K=2.62 tau=9.802467865447825e-08 off=-0.2

*Grain_499:
XU_499 in out fe_tanh Vc=0.3703603018652145 Qo=1.3058573625765125e-13 K=2.62 tau=9.072608644502309e-08 off=-0.2

*Grain_500:
XU_500 in out fe_tanh Vc=0.23447245232061167 Qo=8.2672893569374e-14 K=2.62 tau=9.953029214904018e-08 off=-0.2

*Grain_501:
XU_501 in out fe_tanh Vc=0.4868815859397231 Qo=1.7167010084512317e-13 K=2.62 tau=9.831068834466908e-08 off=-0.2

*Grain_502:
XU_502 in out fe_tanh Vc=0.5173195253436911 Qo=1.824022465616462e-13 K=2.62 tau=8.575937786391419e-08 off=-0.2

*Grain_503:
XU_503 in out fe_tanh Vc=-0.1322794351842998 Qo=4.6640547996892266e-14 K=2.62 tau=1.0162121339157471e-07 off=-0.2

*Grain_504:
XU_504 in out fe_tanh Vc=0.7548061420080543 Qo=2.6613790757139666e-13 K=2.62 tau=1.092558245478408e-07 off=-0.2

*Grain_505:
XU_505 in out fe_tanh Vc=0.7215400451558996 Qo=2.5440857878540306e-13 K=2.62 tau=1.0194715668203179e-07 off=-0.2

*Grain_506:
XU_506 in out fe_tanh Vc=0.18770851999078153 Qo=6.618434848816745e-14 K=2.62 tau=8.814139883656223e-08 off=-0.2

*Grain_507:
XU_507 in out fe_tanh Vc=-0.01196277977442467 Qo=4.217969357579543e-15 K=2.62 tau=1.051169776313394e-07 off=-0.2

*Grain_508:
XU_508 in out fe_tanh Vc=0.41858189973383264 Qo=1.4758824119535805e-13 K=2.62 tau=1.0597038320486302e-07 off=-0.2

*Grain_509:
XU_509 in out fe_tanh Vc=0.12654412459758296 Qo=4.461832868272483e-14 K=2.62 tau=9.318034440384229e-08 off=-0.2

*Grain_510:
XU_510 in out fe_tanh Vc=1.0858136243773848 Qo=3.828481909746146e-13 K=2.62 tau=1.2093691782210417e-07 off=-0.2

*Grain_511:
XU_511 in out fe_tanh Vc=0.7805178449693555 Qo=2.752036245090113e-13 K=2.62 tau=1.0286109239275097e-07 off=-0.2

*Grain_512:
XU_512 in out fe_tanh Vc=0.6808777337382272 Qo=2.4007141076908823e-13 K=2.62 tau=8.837068160437701e-08 off=-0.2

*Grain_513:
XU_513 in out fe_tanh Vc=0.47836592429937047 Qo=1.686675545694395e-13 K=2.62 tau=1.1971729225268535e-07 off=-0.2

*Grain_514:
XU_514 in out fe_tanh Vc=0.7262019068753034 Qo=2.560523096115574e-13 K=2.62 tau=8.822014075306398e-08 off=-0.2

*Grain_515:
XU_515 in out fe_tanh Vc=0.5813190742057203 Qo=2.0496791617098552e-13 K=2.62 tau=1.1174151261877522e-07 off=-0.2

*Grain_516:
XU_516 in out fe_tanh Vc=0.526735589303767 Qo=1.8572226665743695e-13 K=2.62 tau=9.827298053470852e-08 off=-0.2

*Grain_517:
XU_517 in out fe_tanh Vc=0.4545810858253743 Qo=1.6028123284906665e-13 K=2.62 tau=8.491014340320446e-08 off=-0.2

*Grain_518:
XU_518 in out fe_tanh Vc=0.35103793056242927 Qo=1.2377284062572092e-13 K=2.62 tau=1.1072062587618916e-07 off=-0.2

*Grain_519:
XU_519 in out fe_tanh Vc=0.3203309081538937 Qo=1.1294581864387217e-13 K=2.62 tau=1.0477653363206852e-07 off=-0.2

*Grain_520:
XU_520 in out fe_tanh Vc=0.48049390549508153 Qo=1.694178617427107e-13 K=2.62 tau=8.674728486238747e-08 off=-0.2

*Grain_521:
XU_521 in out fe_tanh Vc=-0.1934430627506643 Qo=6.820629707344754e-14 K=2.62 tau=1.1237441496669077e-07 off=-0.2

*Grain_522:
XU_522 in out fe_tanh Vc=0.1416920030901513 Qo=4.9959335415172536e-14 K=2.62 tau=1.1413458555873503e-07 off=-0.2

*Grain_523:
XU_523 in out fe_tanh Vc=-0.3064047880281901 Qo=1.0803559300503108e-13 K=2.62 tau=8.968153554095161e-08 off=-0.2

*Grain_524:
XU_524 in out fe_tanh Vc=0.8453956543855035 Qo=2.980789609495635e-13 K=2.62 tau=1.0307275407064376e-07 off=-0.2

*Grain_525:
XU_525 in out fe_tanh Vc=0.2851152457723637 Qo=1.0052909045585335e-13 K=2.62 tau=8.609489031804692e-08 off=-0.2

*Grain_526:
XU_526 in out fe_tanh Vc=0.1567749375069849 Qo=5.5277443446267315e-14 K=2.62 tau=9.704553426491052e-08 off=-0.2

*Grain_527:
XU_527 in out fe_tanh Vc=0.5276447241347606 Qo=1.8604281948306347e-13 K=2.62 tau=8.118167870391765e-08 off=-0.2

*Grain_528:
XU_528 in out fe_tanh Vc=0.5780822674609816 Qo=2.0382664700753382e-13 K=2.62 tau=1.14346656225066e-07 off=-0.2

*Grain_529:
XU_529 in out fe_tanh Vc=0.4002042353857477 Qo=1.4110844080232334e-13 K=2.62 tau=8.986753368812875e-08 off=-0.2

*Grain_530:
XU_530 in out fe_tanh Vc=0.1465417593036607 Qo=5.166931616262782e-14 K=2.62 tau=1.1415749953935951e-07 off=-0.2

*Grain_531:
XU_531 in out fe_tanh Vc=0.4001000840822592 Qo=1.4107171798246457e-13 K=2.62 tau=1.0293950031057128e-07 off=-0.2

*Grain_532:
XU_532 in out fe_tanh Vc=0.7352570988326286 Qo=2.5924508946065693e-13 K=2.62 tau=8.926602435740144e-08 off=-0.2

*Grain_533:
XU_533 in out fe_tanh Vc=0.591118205351345 Qo=2.0842300233678733e-13 K=2.62 tau=1.1130213732238235e-07 off=-0.2

*Grain_534:
XU_534 in out fe_tanh Vc=0.004685773727148845 Qo=1.6521619866245222e-15 K=2.62 tau=9.552986114697173e-08 off=-0.2

*Grain_535:
XU_535 in out fe_tanh Vc=0.6184064418176096 Qo=2.1804459091464983e-13 K=2.62 tau=1.1391931085449605e-07 off=-0.2

*Grain_536:
XU_536 in out fe_tanh Vc=0.3333168742579979 Qo=1.1752455436738523e-13 K=2.62 tau=1.0505256948150295e-07 off=-0.2

*Grain_537:
XU_537 in out fe_tanh Vc=0.47912229318963045 Qo=1.6893424348809398e-13 K=2.62 tau=1.1602693675787364e-07 off=-0.2

*Grain_538:
XU_538 in out fe_tanh Vc=0.6346405149594654 Qo=2.2376858018405404e-13 K=2.62 tau=1.1010743284640556e-07 off=-0.2

*Grain_539:
XU_539 in out fe_tanh Vc=0.476269169036929 Qo=1.6792825738148746e-13 K=2.62 tau=8.769983141321268e-08 off=-0.2

*Grain_540:
XU_540 in out fe_tanh Vc=0.6404176027595052 Qo=2.2580552977069698e-13 K=2.62 tau=8.358867454093651e-08 off=-0.2

*Grain_541:
XU_541 in out fe_tanh Vc=0.3290421784780201 Qo=1.160173347952697e-13 K=2.62 tau=9.297539779627079e-08 off=-0.2

*Grain_542:
XU_542 in out fe_tanh Vc=0.27944399040867984 Qo=9.852945644151092e-14 K=2.62 tau=1.1243165027173678e-07 off=-0.2

*Grain_543:
XU_543 in out fe_tanh Vc=0.5363324384819942 Qo=1.8910603000729113e-13 K=2.62 tau=1.081745586416968e-07 off=-0.2

*Grain_544:
XU_544 in out fe_tanh Vc=0.4208372708532601 Qo=1.4838346491853088e-13 K=2.62 tau=8.913265985155215e-08 off=-0.2

*Grain_545:
XU_545 in out fe_tanh Vc=0.3267328482718872 Qo=1.1520308557981342e-13 K=2.62 tau=9.663815451406869e-08 off=-0.2

*Grain_546:
XU_546 in out fe_tanh Vc=0.9035931340209291 Qo=3.18598872744261e-13 K=2.62 tau=9.390569995697197e-08 off=-0.2

*Grain_547:
XU_547 in out fe_tanh Vc=0.02866409633737438 Qo=1.0106704486212766e-14 K=2.62 tau=8.930958726304875e-08 off=-0.2

*Grain_548:
XU_548 in out fe_tanh Vc=0.8535284719235323 Qo=3.0094651981238986e-13 K=2.62 tau=9.14003402785387e-08 off=-0.2

*Grain_549:
XU_549 in out fe_tanh Vc=1.0775103228114404 Qo=3.7992052096544404e-13 K=2.62 tau=1.0041055982812095e-07 off=-0.2

*Grain_550:
XU_550 in out fe_tanh Vc=0.19750799724706763 Qo=6.963955668949877e-14 K=2.62 tau=1.0000018163599317e-07 off=-0.2

*Grain_551:
XU_551 in out fe_tanh Vc=0.21518709500369432 Qo=7.587304873843946e-14 K=2.62 tau=1.0800172217985703e-07 off=-0.2

*Grain_552:
XU_552 in out fe_tanh Vc=0.8268535148883074 Qo=2.915411680872102e-13 K=2.62 tau=1.0853953921772501e-07 off=-0.2

*Grain_553:
XU_553 in out fe_tanh Vc=0.22772335470794652 Qo=8.029322199986171e-14 K=2.62 tau=1.0318446224995569e-07 off=-0.2

*Grain_554:
XU_554 in out fe_tanh Vc=0.4923895601791405 Qo=1.736121633926482e-13 K=2.62 tau=1.073275035846719e-07 off=-0.2

*Grain_555:
XU_555 in out fe_tanh Vc=0.28202325248973725 Qo=9.943888122640296e-14 K=2.62 tau=8.740220756988443e-08 off=-0.2

*Grain_556:
XU_556 in out fe_tanh Vc=0.31904527263728155 Qo=1.1249251503749137e-13 K=2.62 tau=9.190175012891577e-08 off=-0.2

*Grain_557:
XU_557 in out fe_tanh Vc=-0.06754611785244918 Qo=2.3816158175392756e-14 K=2.62 tau=8.885051858217613e-08 off=-0.2

*Grain_558:
XU_558 in out fe_tanh Vc=-0.023899839151030666 Qo=8.42686993249238e-15 K=2.62 tau=8.751780218564785e-08 off=-0.2

*Grain_559:
XU_559 in out fe_tanh Vc=0.3123158573559896 Qo=1.1011978328231851e-13 K=2.62 tau=1.0052514878865054e-07 off=-0.2

*Grain_560:
XU_560 in out fe_tanh Vc=0.5769139807286805 Qo=2.0341471953493686e-13 K=2.62 tau=9.529528118784894e-08 off=-0.2

*Grain_561:
XU_561 in out fe_tanh Vc=0.15645581613553783 Qo=5.516492409946882e-14 K=2.62 tau=8.596554146173647e-08 off=-0.2

*Grain_562:
XU_562 in out fe_tanh Vc=0.4956844646654436 Qo=1.7477391730114112e-13 K=2.62 tau=9.353569778017117e-08 off=-0.2

*Grain_563:
XU_563 in out fe_tanh Vc=0.6501769178576362 Qo=2.292465771535875e-13 K=2.62 tau=9.694516064332975e-08 off=-0.2

*Grain_564:
XU_564 in out fe_tanh Vc=0.23854556565502796 Qo=8.410903697069668e-14 K=2.62 tau=9.751168960203018e-08 off=-0.2

*Grain_565:
XU_565 in out fe_tanh Vc=0.29769912960844047 Qo=1.0496605556101972e-13 K=2.62 tau=8.322069224240833e-08 off=-0.2

*Grain_566:
XU_566 in out fe_tanh Vc=0.12111215014240939 Qo=4.270306298067951e-14 K=2.62 tau=1.0017300911464129e-07 off=-0.2

*Grain_567:
XU_567 in out fe_tanh Vc=0.5288814470892967 Qo=1.8647887695669522e-13 K=2.62 tau=9.985296460616523e-08 off=-0.2

*Grain_568:
XU_568 in out fe_tanh Vc=0.5689623787602155 Qo=2.0061105566424025e-13 K=2.62 tau=9.341774751361589e-08 off=-0.2

*Grain_569:
XU_569 in out fe_tanh Vc=0.8043888299354515 Qo=2.83620320713475e-13 K=2.62 tau=9.472316814467621e-08 off=-0.2

*Grain_570:
XU_570 in out fe_tanh Vc=0.5528595610579377 Qo=1.9493334589112326e-13 K=2.62 tau=8.979798304477145e-08 off=-0.2

*Grain_571:
XU_571 in out fe_tanh Vc=0.5118801453195229 Qo=1.8048436972208237e-13 K=2.62 tau=1.0780121147665401e-07 off=-0.2

*Grain_572:
XU_572 in out fe_tanh Vc=0.7420396364028654 Qo=2.616365516606929e-13 K=2.62 tau=1.0735119954891635e-07 off=-0.2

*Grain_573:
XU_573 in out fe_tanh Vc=0.48082570260701935 Qo=1.6953485044245084e-13 K=2.62 tau=9.438334895582324e-08 off=-0.2

*Grain_574:
XU_574 in out fe_tanh Vc=0.2933276763823154 Qo=1.0342472017713946e-13 K=2.62 tau=1.048083427736363e-07 off=-0.2

*Grain_575:
XU_575 in out fe_tanh Vc=0.4014155451983165 Qo=1.4153553782895873e-13 K=2.62 tau=1.0460193095165477e-07 off=-0.2

*Grain_576:
XU_576 in out fe_tanh Vc=0.8223057909755564 Qo=2.8993768123278153e-13 K=2.62 tau=1.0854616571391616e-07 off=-0.2

*Grain_577:
XU_577 in out fe_tanh Vc=-0.0542212512773233 Qo=1.9117929171137774e-14 K=2.62 tau=9.392799974264955e-08 off=-0.2

*Grain_578:
XU_578 in out fe_tanh Vc=0.706427136387179 Qo=2.490799020654118e-13 K=2.62 tau=1.1123771259376522e-07 off=-0.2

*Grain_579:
XU_579 in out fe_tanh Vc=0.4051723533034259 Qo=1.4286015483006203e-13 K=2.62 tau=1.0621831888090526e-07 off=-0.2

*Grain_580:
XU_580 in out fe_tanh Vc=0.6759986200521636 Qo=2.383510788388824e-13 K=2.62 tau=1.1927776336198525e-07 off=-0.2

*Grain_581:
XU_581 in out fe_tanh Vc=0.9835970964883294 Qo=3.468075557205944e-13 K=2.62 tau=1.1479565523485088e-07 off=-0.2

*Grain_582:
XU_582 in out fe_tanh Vc=0.49371923449627464 Qo=1.7408099468696182e-13 K=2.62 tau=1.0881023743939635e-07 off=-0.2

*Grain_583:
XU_583 in out fe_tanh Vc=0.26783580928059203 Qo=9.443651540115291e-14 K=2.62 tau=1.117670626299416e-07 off=-0.2

*Grain_584:
XU_584 in out fe_tanh Vc=0.6108343196425959 Qo=2.153747282315351e-13 K=2.62 tau=1.1118510187211033e-07 off=-0.2

*Grain_585:
XU_585 in out fe_tanh Vc=0.9476401003910491 Qo=3.341294398822352e-13 K=2.62 tau=1.0494431289234571e-07 off=-0.2

*Grain_586:
XU_586 in out fe_tanh Vc=0.6549905164021576 Qo=2.3094380902973454e-13 K=2.62 tau=9.061921224765627e-08 off=-0.2

*Grain_587:
XU_587 in out fe_tanh Vc=0.010472598672029987 Qo=3.692544803615691e-15 K=2.62 tau=1.0468359397504554e-07 off=-0.2

*Grain_588:
XU_588 in out fe_tanh Vc=0.46110018911914796 Qo=1.6257981047488065e-13 K=2.62 tau=9.240150564199147e-08 off=-0.2

*Grain_589:
XU_589 in out fe_tanh Vc=0.2787022323988338 Qo=9.82679191888601e-14 K=2.62 tau=8.95143926209609e-08 off=-0.2

*Grain_590:
XU_590 in out fe_tanh Vc=0.25891051395129777 Qo=9.128953594351915e-14 K=2.62 tau=9.495206360711114e-08 off=-0.2

*Grain_591:
XU_591 in out fe_tanh Vc=0.6425919489882925 Qo=2.2657218484073354e-13 K=2.62 tau=6.987973955122868e-08 off=-0.2

*Grain_592:
XU_592 in out fe_tanh Vc=0.5374692769639919 Qo=1.895068691075674e-13 K=2.62 tau=1.0840124467038753e-07 off=-0.2

*Grain_593:
XU_593 in out fe_tanh Vc=0.8465950179118301 Qo=2.9850184582231356e-13 K=2.62 tau=9.778192554064522e-08 off=-0.2

*Grain_594:
XU_594 in out fe_tanh Vc=0.36918171422321744 Qo=1.3017017677625098e-13 K=2.62 tau=1.0377559140749891e-07 off=-0.2

*Grain_595:
XU_595 in out fe_tanh Vc=0.36688079461159817 Qo=1.2935889306133943e-13 K=2.62 tau=1.0008292813308527e-07 off=-0.2

*Grain_596:
XU_596 in out fe_tanh Vc=0.7444425975026583 Qo=2.6248381429341737e-13 K=2.62 tau=9.992585329578957e-08 off=-0.2

*Grain_597:
XU_597 in out fe_tanh Vc=0.9623603604078794 Qo=3.393196721574574e-13 K=2.62 tau=9.322588449244285e-08 off=-0.2

*Grain_598:
XU_598 in out fe_tanh Vc=0.15436530560260248 Qo=5.4427828747394376e-14 K=2.62 tau=1.0424619168206146e-07 off=-0.2

*Grain_599:
XU_599 in out fe_tanh Vc=0.6416515564428342 Qo=2.262406108240222e-13 K=2.62 tau=1.0682940074848911e-07 off=-0.2

*Grain_600:
XU_600 in out fe_tanh Vc=0.39633678529657834 Qo=1.397448124253336e-13 K=2.62 tau=1.1344327776141547e-07 off=-0.2

*Grain_601:
XU_601 in out fe_tanh Vc=0.38542257766983506 Qo=1.3589656024649767e-13 K=2.62 tau=9.693284475004099e-08 off=-0.2

*Grain_602:
XU_602 in out fe_tanh Vc=0.5223944394436254 Qo=1.841916159698865e-13 K=2.62 tau=8.127661708322425e-08 off=-0.2

*Grain_603:
XU_603 in out fe_tanh Vc=0.5026972820866628 Qo=1.7724657412094162e-13 K=2.62 tau=9.350592775902412e-08 off=-0.2

*Grain_604:
XU_604 in out fe_tanh Vc=0.2305408225498761 Qo=8.128663600959143e-14 K=2.62 tau=9.984475815187348e-08 off=-0.2

*Grain_605:
XU_605 in out fe_tanh Vc=0.097989053885297 Qo=3.4550065658654247e-14 K=2.62 tau=9.524278240545443e-08 off=-0.2

*Grain_606:
XU_606 in out fe_tanh Vc=0.3684203273716115 Qo=1.299017185692209e-13 K=2.62 tau=1.0162554373763045e-07 off=-0.2

*Grain_607:
XU_607 in out fe_tanh Vc=0.6517865084384397 Qo=2.298141044236784e-13 K=2.62 tau=8.721772049809766e-08 off=-0.2

*Grain_608:
XU_608 in out fe_tanh Vc=0.3454709962513757 Qo=1.218099892832693e-13 K=2.62 tau=1.1233677876637476e-07 off=-0.2

*Grain_609:
XU_609 in out fe_tanh Vc=0.7244060819665215 Qo=2.5541911777992195e-13 K=2.62 tau=1.0378951399451226e-07 off=-0.2

*Grain_610:
XU_610 in out fe_tanh Vc=0.4169629845917266 Qo=1.4701742616819154e-13 K=2.62 tau=9.202575347422794e-08 off=-0.2

*Grain_611:
XU_611 in out fe_tanh Vc=0.18704341421303466 Qo=6.59498381282858e-14 K=2.62 tau=9.048566696265743e-08 off=-0.2

*Grain_612:
XU_612 in out fe_tanh Vc=0.4029766121803692 Qo=1.4208595611129679e-13 K=2.62 tau=9.090715260082878e-08 off=-0.2

*Grain_613:
XU_613 in out fe_tanh Vc=0.28503694321904854 Qo=1.0050148167455574e-13 K=2.62 tau=9.926934115533897e-08 off=-0.2

*Grain_614:
XU_614 in out fe_tanh Vc=0.9446782915948754 Qo=3.3308513254056045e-13 K=2.62 tau=9.73899578872376e-08 off=-0.2

*Grain_615:
XU_615 in out fe_tanh Vc=0.7026724608098004 Qo=2.477560369745494e-13 K=2.62 tau=9.669745309417345e-08 off=-0.2

*Grain_616:
XU_616 in out fe_tanh Vc=0.3384798138906608 Qo=1.19344960792668e-13 K=2.62 tau=1.0020440201417908e-07 off=-0.2

*Grain_617:
XU_617 in out fe_tanh Vc=0.3863562862275162 Qo=1.3622577754878629e-13 K=2.62 tau=1.0398419973803146e-07 off=-0.2

*Grain_618:
XU_618 in out fe_tanh Vc=0.6950005506369707 Qo=2.4505098993420515e-13 K=2.62 tau=7.821094819052147e-08 off=-0.2

*Grain_619:
XU_619 in out fe_tanh Vc=0.5099140936278124 Qo=1.797911574463886e-13 K=2.62 tau=9.144854848045013e-08 off=-0.2

*Grain_620:
XU_620 in out fe_tanh Vc=-0.11655048555199682 Qo=4.1094660767754785e-14 K=2.62 tau=9.700525762755328e-08 off=-0.2

*Grain_621:
XU_621 in out fe_tanh Vc=0.6910096622060962 Qo=2.436438382998554e-13 K=2.62 tau=1.047578286510961e-07 off=-0.2

*Grain_622:
XU_622 in out fe_tanh Vc=0.4027952104868105 Qo=1.42021995493508e-13 K=2.62 tau=1.073423046792884e-07 off=-0.2

*Grain_623:
XU_623 in out fe_tanh Vc=1.1090729774728012 Qo=3.910492312414708e-13 K=2.62 tau=9.352017457042885e-08 off=-0.2

*Grain_624:
XU_624 in out fe_tanh Vc=-0.0014464535188143945 Qo=5.100065983464654e-16 K=2.62 tau=1.0501839801464848e-07 off=-0.2

*Grain_625:
XU_625 in out fe_tanh Vc=0.840400646052901 Qo=2.963177656015714e-13 K=2.62 tau=1.0551786558020826e-07 off=-0.2

*Grain_626:
XU_626 in out fe_tanh Vc=0.917743780978292 Qo=3.2358826453961014e-13 K=2.62 tau=1.0946411597027255e-07 off=-0.2

*Grain_627:
XU_627 in out fe_tanh Vc=0.2827729273530442 Qo=9.970320989091091e-14 K=2.62 tau=9.969434277021671e-08 off=-0.2

*Grain_628:
XU_628 in out fe_tanh Vc=0.4092060165088632 Qo=1.4428238846807522e-13 K=2.62 tau=9.467998366477285e-08 off=-0.2

*Grain_629:
XU_629 in out fe_tanh Vc=1.1147493339732295 Qo=3.9305066387109186e-13 K=2.62 tau=1.0335018034308475e-07 off=-0.2

*Grain_630:
XU_630 in out fe_tanh Vc=0.14951911906880916 Qo=5.271910663714071e-14 K=2.62 tau=1.0078335417287834e-07 off=-0.2

*Grain_631:
XU_631 in out fe_tanh Vc=0.43363685620398396 Qo=1.5289648445220977e-13 K=2.62 tau=1.0743742608614269e-07 off=-0.2

*Grain_632:
XU_632 in out fe_tanh Vc=0.5682134962339047 Qo=2.0034700637068402e-13 K=2.62 tau=1.0441484261920552e-07 off=-0.2

*Grain_633:
XU_633 in out fe_tanh Vc=0.16720732744330313 Qo=5.895581100861156e-14 K=2.62 tau=9.390359332243609e-08 off=-0.2

*Grain_634:
XU_634 in out fe_tanh Vc=0.7373169643292325 Qo=2.59971379646487e-13 K=2.62 tau=9.641304956423783e-08 off=-0.2

*Grain_635:
XU_635 in out fe_tanh Vc=0.2260732077118108 Qo=7.971139489976891e-14 K=2.62 tau=9.298329207872579e-08 off=-0.2

*Grain_636:
XU_636 in out fe_tanh Vc=0.09101591630709022 Qo=3.20913995972808e-14 K=2.62 tau=1.0114953676084189e-07 off=-0.2

*Grain_637:
XU_637 in out fe_tanh Vc=0.37836184713727355 Qo=1.3340700969135478e-13 K=2.62 tau=9.641226846937362e-08 off=-0.2

*Grain_638:
XU_638 in out fe_tanh Vc=0.12592480195910688 Qo=4.4399961049047224e-14 K=2.62 tau=1.0348520819577384e-07 off=-0.2

*Grain_639:
XU_639 in out fe_tanh Vc=0.0360160538004638 Qo=1.2698939057297712e-14 K=2.62 tau=1.0790061769874062e-07 off=-0.2

*Grain_640:
XU_640 in out fe_tanh Vc=0.32042516983818226 Qo=1.1297905447228497e-13 K=2.62 tau=1.0661740897522522e-07 off=-0.2

*Grain_641:
XU_641 in out fe_tanh Vc=0.3472471951773258 Qo=1.2243626116855808e-13 K=2.62 tau=1.1063012135159052e-07 off=-0.2

*Grain_642:
XU_642 in out fe_tanh Vc=0.6327294683193457 Qo=2.2309476219852504e-13 K=2.62 tau=1.0801339771775188e-07 off=-0.2

*Grain_643:
XU_643 in out fe_tanh Vc=0.38497226524252753 Qo=1.3573778410453597e-13 K=2.62 tau=8.402163014365919e-08 off=-0.2

*Grain_644:
XU_644 in out fe_tanh Vc=0.7005833101443245 Qo=2.4701942109960174e-13 K=2.62 tau=9.063002658593455e-08 off=-0.2

*Grain_645:
XU_645 in out fe_tanh Vc=0.7965228204702322 Qo=2.808468359953446e-13 K=2.62 tau=1.0131744377859137e-07 off=-0.2

*Grain_646:
XU_646 in out fe_tanh Vc=0.27614344141613567 Qo=9.736571233050551e-14 K=2.62 tau=1.1090283120918054e-07 off=-0.2

*Grain_647:
XU_647 in out fe_tanh Vc=-0.05911773756758326 Qo=2.084438652649924e-14 K=2.62 tau=1.0724166372012618e-07 off=-0.2

*Grain_648:
XU_648 in out fe_tanh Vc=0.5789407643808009 Qo=2.0412934535772128e-13 K=2.62 tau=9.050617427528985e-08 off=-0.2

*Grain_649:
XU_649 in out fe_tanh Vc=0.3183853343765358 Qo=1.1225982669797425e-13 K=2.62 tau=1.1940443973812807e-07 off=-0.2

*Grain_650:
XU_650 in out fe_tanh Vc=0.1591921769536146 Qo=5.6129740496624656e-14 K=2.62 tau=9.168747008269255e-08 off=-0.2

*Grain_651:
XU_651 in out fe_tanh Vc=0.55374522178055 Qo=1.952456219556862e-13 K=2.62 tau=1.1528131649004071e-07 off=-0.2

*Grain_652:
XU_652 in out fe_tanh Vc=0.6446914160469677 Qo=2.2731243818382958e-13 K=2.62 tau=9.015816676438711e-08 off=-0.2

*Grain_653:
XU_653 in out fe_tanh Vc=0.2955797376892173 Qo=1.0421877688996227e-13 K=2.62 tau=9.648371903000647e-08 off=-0.2

*Grain_654:
XU_654 in out fe_tanh Vc=0.05044928817173999 Qo=1.7787968652154957e-14 K=2.62 tau=1.0572874037062859e-07 off=-0.2

*Grain_655:
XU_655 in out fe_tanh Vc=0.8344091317723205 Qo=2.9420521115205974e-13 K=2.62 tau=1.0341563993817188e-07 off=-0.2

*Grain_656:
XU_656 in out fe_tanh Vc=0.44330365519515424 Qo=1.5630491148167065e-13 K=2.62 tau=9.043854333119065e-08 off=-0.2

*Grain_657:
XU_657 in out fe_tanh Vc=0.3490515306290218 Qo=1.2307245374165207e-13 K=2.62 tau=1.064505920327449e-07 off=-0.2

*Grain_658:
XU_658 in out fe_tanh Vc=0.8230661927582101 Qo=2.902057921132927e-13 K=2.62 tau=1.050372271002234e-07 off=-0.2

*Grain_659:
XU_659 in out fe_tanh Vc=0.361994126659185 Qo=1.2763589756425514e-13 K=2.62 tau=9.983869038401639e-08 off=-0.2

*Grain_660:
XU_660 in out fe_tanh Vc=0.6402077640101441 Qo=2.2573154250088783e-13 K=2.62 tau=1.0243768423287621e-07 off=-0.2

*Grain_661:
XU_661 in out fe_tanh Vc=-0.03866174635638342 Qo=1.3631786634606053e-14 K=2.62 tau=1.0369414400891322e-07 off=-0.2

*Grain_662:
XU_662 in out fe_tanh Vc=0.41774089028323985 Qo=1.4729170877071046e-13 K=2.62 tau=1.0116045651215319e-07 off=-0.2

*Grain_663:
XU_663 in out fe_tanh Vc=0.27192728010562606 Qo=9.587913148979141e-14 K=2.62 tau=9.168395024851822e-08 off=-0.2

*Grain_664:
XU_664 in out fe_tanh Vc=0.4735679648837188 Qo=1.6697583691052252e-13 K=2.62 tau=1.0987012802294467e-07 off=-0.2

*Grain_665:
XU_665 in out fe_tanh Vc=0.7809737870959154 Qo=2.753643856326735e-13 K=2.62 tau=1.0992715924529682e-07 off=-0.2

*Grain_666:
XU_666 in out fe_tanh Vc=-0.015777223755437775 Qo=5.5629082540151575e-15 K=2.62 tau=1.0677707714056269e-07 off=-0.2

*Grain_667:
XU_667 in out fe_tanh Vc=0.5801897017645632 Qo=2.0456970953006086e-13 K=2.62 tau=8.704625796189015e-08 off=-0.2

*Grain_668:
XU_668 in out fe_tanh Vc=0.2849566007350033 Qo=1.0047315363189302e-13 K=2.62 tau=1.0373575556827398e-07 off=-0.2

*Grain_669:
XU_669 in out fe_tanh Vc=0.4347067199416999 Qo=1.5327370885553106e-13 K=2.62 tau=9.064279272442432e-08 off=-0.2

*Grain_670:
XU_670 in out fe_tanh Vc=0.2665805681597819 Qo=9.39939285874033e-14 K=2.62 tau=1.2483323849563228e-07 off=-0.2

*Grain_671:
XU_671 in out fe_tanh Vc=0.019807130466933276 Qo=6.983817385798424e-15 K=2.62 tau=8.890132637876362e-08 off=-0.2

*Grain_672:
XU_672 in out fe_tanh Vc=0.1509511131545444 Qo=5.322401496846179e-14 K=2.62 tau=1.0553627302975135e-07 off=-0.2

*Grain_673:
XU_673 in out fe_tanh Vc=0.9771361527599844 Qo=3.445294846383642e-13 K=2.62 tau=1.0307115629070717e-07 off=-0.2

*Grain_674:
XU_674 in out fe_tanh Vc=-0.051873356523848 Qo=1.829008244055154e-14 K=2.62 tau=7.625381509773376e-08 off=-0.2

*Grain_675:
XU_675 in out fe_tanh Vc=-0.040690998213741225 Qo=1.4347282724523685e-14 K=2.62 tau=9.785812770376124e-08 off=-0.2

*Grain_676:
XU_676 in out fe_tanh Vc=0.7910332142346144 Qo=2.789112498419895e-13 K=2.62 tau=9.622026013561653e-08 off=-0.2

*Grain_677:
XU_677 in out fe_tanh Vc=0.4436063397756938 Qo=1.5641163536272524e-13 K=2.62 tau=9.653969618714437e-08 off=-0.2

*Grain_678:
XU_678 in out fe_tanh Vc=0.5903393146797475 Qo=2.081483724390836e-13 K=2.62 tau=9.407844312036506e-08 off=-0.2

*Grain_679:
XU_679 in out fe_tanh Vc=0.9033808112088386 Qo=3.1852400961610854e-13 K=2.62 tau=1.277522530176775e-07 off=-0.2

*Grain_680:
XU_680 in out fe_tanh Vc=0.5188350954157422 Qo=1.829366230396654e-13 K=2.62 tau=8.145356004932649e-08 off=-0.2

*Grain_681:
XU_681 in out fe_tanh Vc=1.0706164587323288 Qo=3.774898060321827e-13 K=2.62 tau=8.953722788582031e-08 off=-0.2

*Grain_682:
XU_682 in out fe_tanh Vc=0.724433022052541 Qo=2.554286166137602e-13 K=2.62 tau=1.0689292393308495e-07 off=-0.2

*Grain_683:
XU_683 in out fe_tanh Vc=0.2726016217774251 Qo=9.611689834346769e-14 K=2.62 tau=9.454779830827259e-08 off=-0.2

*Grain_684:
XU_684 in out fe_tanh Vc=0.05618294700892734 Qo=1.980960557418335e-14 K=2.62 tau=1.1413905330666704e-07 off=-0.2

*Grain_685:
XU_685 in out fe_tanh Vc=0.41591857702124013 Qo=1.4664917738218998e-13 K=2.62 tau=1.0616559864760392e-07 off=-0.2

*Grain_686:
XU_686 in out fe_tanh Vc=-0.002474192296872235 Qo=8.723781169388234e-16 K=2.62 tau=1.0014744335477048e-07 off=-0.2

*Grain_687:
XU_687 in out fe_tanh Vc=0.2503426816012191 Qo=8.826859474131028e-14 K=2.62 tau=9.5680388455628e-08 off=-0.2

*Grain_688:
XU_688 in out fe_tanh Vc=0.2823136995213913 Qo=9.954129025696423e-14 K=2.62 tau=1.0637559325383278e-07 off=-0.2

*Grain_689:
XU_689 in out fe_tanh Vc=0.614972625307287 Qo=2.1683385786654538e-13 K=2.62 tau=1.1207015226129012e-07 off=-0.2

*Grain_690:
XU_690 in out fe_tanh Vc=0.610990916906281 Qo=2.1542994302877784e-13 K=2.62 tau=1.0429070467253712e-07 off=-0.2

*Grain_691:
XU_691 in out fe_tanh Vc=0.5958742273654217 Qo=2.1009993324228119e-13 K=2.62 tau=1.0747700667857444e-07 off=-0.2

*Grain_692:
XU_692 in out fe_tanh Vc=0.47287021825032166 Qo=1.6672981767632116e-13 K=2.62 tau=1.0303836923629264e-07 off=-0.2

*Grain_693:
XU_693 in out fe_tanh Vc=0.5843326432870442 Qo=2.060304737271439e-13 K=2.62 tau=7.323190223486317e-08 off=-0.2

*Grain_694:
XU_694 in out fe_tanh Vc=0.6807896300396887 Qo=2.40040346191479e-13 K=2.62 tau=9.438228266079737e-08 off=-0.2

*Grain_695:
XU_695 in out fe_tanh Vc=0.6140327682265436 Qo=2.1650247264991246e-13 K=2.62 tau=9.454730125764727e-08 off=-0.2

*Grain_696:
XU_696 in out fe_tanh Vc=0.36460009005549593 Qo=1.2855473699454484e-13 K=2.62 tau=9.396119230048093e-08 off=-0.2

*Grain_697:
XU_697 in out fe_tanh Vc=0.829726338854346 Qo=2.925541001721406e-13 K=2.62 tau=8.957315615098377e-08 off=-0.2

*Grain_698:
XU_698 in out fe_tanh Vc=0.7829041695360553 Qo=2.7604502124868036e-13 K=2.62 tau=1.1156296725920179e-07 off=-0.2

*Grain_699:
XU_699 in out fe_tanh Vc=-0.019744011849928078 Qo=6.961562324897787e-15 K=2.62 tau=9.703013893061202e-08 off=-0.2

*Grain_700:
XU_700 in out fe_tanh Vc=0.06578856406144046 Qo=2.319646039824053e-14 K=2.62 tau=1.0089830820775479e-07 off=-0.2

*Grain_701:
XU_701 in out fe_tanh Vc=0.7158688333184304 Qo=2.524089601180154e-13 K=2.62 tau=9.940936132247464e-08 off=-0.2

*Grain_702:
XU_702 in out fe_tanh Vc=0.43221849767054393 Qo=1.5239638389490437e-13 K=2.62 tau=9.441910817089733e-08 off=-0.2

*Grain_703:
XU_703 in out fe_tanh Vc=0.3309978506602319 Qo=1.1670688734857138e-13 K=2.62 tau=9.268488554544654e-08 off=-0.2

*Grain_704:
XU_704 in out fe_tanh Vc=0.17912705911608884 Qo=6.315860198984055e-14 K=2.62 tau=8.847436157105512e-08 off=-0.2

*Grain_705:
XU_705 in out fe_tanh Vc=0.6968764262759752 Qo=2.4571240693870995e-13 K=2.62 tau=8.888114095105015e-08 off=-0.2

*Grain_706:
XU_706 in out fe_tanh Vc=0.4682135835745047 Qo=1.6508792985907404e-13 K=2.62 tau=1.0060573246459854e-07 off=-0.2

*Grain_707:
XU_707 in out fe_tanh Vc=0.30135694226737975 Qo=1.0625576765152875e-13 K=2.62 tau=9.873157774550647e-08 off=-0.2

*Grain_708:
XU_708 in out fe_tanh Vc=0.49414073165488753 Qo=1.7422961082241366e-13 K=2.62 tau=1.0637499578406196e-07 off=-0.2

*Grain_709:
XU_709 in out fe_tanh Vc=0.8244762775170212 Qo=2.9070297541152333e-13 K=2.62 tau=9.971007710239884e-08 off=-0.2

*Grain_710:
XU_710 in out fe_tanh Vc=0.38534197033302914 Qo=1.3586813881911585e-13 K=2.62 tau=9.308369029072813e-08 off=-0.2

*Grain_711:
XU_711 in out fe_tanh Vc=0.3692242237097856 Qo=1.3018516524173574e-13 K=2.62 tau=1.0422801457862982e-07 off=-0.2

*Grain_712:
XU_712 in out fe_tanh Vc=0.17915659415015295 Qo=6.31690157791944e-14 K=2.62 tau=8.6334223495619e-08 off=-0.2

*Grain_713:
XU_713 in out fe_tanh Vc=0.2665709366789174 Qo=9.399053261323002e-14 K=2.62 tau=1.0676132844378034e-07 off=-0.2

*Grain_714:
XU_714 in out fe_tanh Vc=1.1032360103845524 Qo=3.8899116875234357e-13 K=2.62 tau=8.582724735706966e-08 off=-0.2

*Grain_715:
XU_715 in out fe_tanh Vc=0.10841897128953765 Qo=3.8227561428260054e-14 K=2.62 tau=1.0165962702267794e-07 off=-0.2

*Grain_716:
XU_716 in out fe_tanh Vc=0.6732274622476541 Qo=2.373739933349406e-13 K=2.62 tau=1.0468461004844468e-07 off=-0.2

*Grain_717:
XU_717 in out fe_tanh Vc=0.7100194200163626 Qo=2.5034650920500196e-13 K=2.62 tau=9.917828173075613e-08 off=-0.2

*Grain_718:
XU_718 in out fe_tanh Vc=0.9363690744531684 Qo=3.301553767521839e-13 K=2.62 tau=1.025311493253972e-07 off=-0.2

*Grain_719:
XU_719 in out fe_tanh Vc=0.4017994399731081 Qo=1.4167089569954894e-13 K=2.62 tau=1.0247047152756983e-07 off=-0.2

*Grain_720:
XU_720 in out fe_tanh Vc=0.029737574033646297 Qo=1.0485203139059344e-14 K=2.62 tau=9.367184724643665e-08 off=-0.2

*Grain_721:
XU_721 in out fe_tanh Vc=0.3188886900633974 Qo=1.1243730541974129e-13 K=2.62 tau=1.1164578537907136e-07 off=-0.2

*Grain_722:
XU_722 in out fe_tanh Vc=0.5629722105457509 Qo=1.9849897582562483e-13 K=2.62 tau=8.99634240366533e-08 off=-0.2

*Grain_723:
XU_723 in out fe_tanh Vc=0.14000876142426255 Qo=4.936583942995857e-14 K=2.62 tau=9.739940834084415e-08 off=-0.2

*Grain_724:
XU_724 in out fe_tanh Vc=0.4832738709322751 Qo=1.703980527393118e-13 K=2.62 tau=1.1179922709623156e-07 off=-0.2

*Grain_725:
XU_725 in out fe_tanh Vc=0.5080937534852537 Qo=1.7914932176216912e-13 K=2.62 tau=1.0948148153736457e-07 off=-0.2

*Grain_726:
XU_726 in out fe_tanh Vc=0.5847981394335173 Qo=2.0619460351293939e-13 K=2.62 tau=1.1220990842648786e-07 off=-0.2

*Grain_727:
XU_727 in out fe_tanh Vc=0.31257974259751886 Qo=1.1021282686279699e-13 K=2.62 tau=1.0646968688100786e-07 off=-0.2

*Grain_728:
XU_728 in out fe_tanh Vc=0.2179550096609305 Qo=7.684899073760402e-14 K=2.62 tau=9.083199232711735e-08 off=-0.2

*Grain_729:
XU_729 in out fe_tanh Vc=0.3446610544459265 Qo=1.215244110329607e-13 K=2.62 tau=1.1080383708295262e-07 off=-0.2

*Grain_730:
XU_730 in out fe_tanh Vc=0.23948655473965763 Qo=8.444082132179459e-14 K=2.62 tau=8.870701234218705e-08 off=-0.2

*Grain_731:
XU_731 in out fe_tanh Vc=0.5974813310617948 Qo=2.1066658365912216e-13 K=2.62 tau=9.36404216521449e-08 off=-0.2

*Grain_732:
XU_732 in out fe_tanh Vc=0.4252070746635115 Qo=1.499242187330983e-13 K=2.62 tau=9.089873357992665e-08 off=-0.2

*Grain_733:
XU_733 in out fe_tanh Vc=0.32054143585482336 Qo=1.1302004883185419e-13 K=2.62 tau=9.372058326412251e-08 off=-0.2

*Grain_734:
XU_734 in out fe_tanh Vc=0.2659882936951189 Qo=9.378509789835507e-14 K=2.62 tau=9.384232693778173e-08 off=-0.2

*Grain_735:
XU_735 in out fe_tanh Vc=0.4379880773396341 Qo=1.54430686181599e-13 K=2.62 tau=8.498530049942736e-08 off=-0.2

*Grain_736:
XU_736 in out fe_tanh Vc=0.6106114676197752 Qo=2.1529615259767264e-13 K=2.62 tau=9.228809139400271e-08 off=-0.2

*Grain_737:
XU_737 in out fe_tanh Vc=0.36260958406798494 Qo=1.2785290235245356e-13 K=2.62 tau=1.0461173869277423e-07 off=-0.2

*Grain_738:
XU_738 in out fe_tanh Vc=-0.04918061011266733 Qo=1.7340644093924568e-14 K=2.62 tau=8.873462937679094e-08 off=-0.2

*Grain_739:
XU_739 in out fe_tanh Vc=0.21775191116244233 Qo=7.677738002008293e-14 K=2.62 tau=1.0848439590000983e-07 off=-0.2

*Grain_740:
XU_740 in out fe_tanh Vc=0.4095537697817023 Qo=1.4440500316770962e-13 K=2.62 tau=1.1064940124620044e-07 off=-0.2

*Grain_741:
XU_741 in out fe_tanh Vc=0.30763160292488373 Qo=1.084681569859161e-13 K=2.62 tau=9.730848854205639e-08 off=-0.2

*Grain_742:
XU_742 in out fe_tanh Vc=0.27363749746750266 Qo=9.648213886460057e-14 K=2.62 tau=9.91189065554463e-08 off=-0.2

*Grain_743:
XU_743 in out fe_tanh Vc=0.0563885729229292 Qo=1.9882107435852525e-14 K=2.62 tau=1.0572673440440834e-07 off=-0.2

*Grain_744:
XU_744 in out fe_tanh Vc=0.24954546588901586 Qo=8.798750359787527e-14 K=2.62 tau=9.956428371308312e-08 off=-0.2

*Grain_745:
XU_745 in out fe_tanh Vc=0.3768443186273217 Qo=1.3287194268561465e-13 K=2.62 tau=1.0219340398818464e-07 off=-0.2

*Grain_746:
XU_746 in out fe_tanh Vc=0.7159709392911826 Qo=2.52444961772515e-13 K=2.62 tau=1.0595557140001593e-07 off=-0.2

*Grain_747:
XU_747 in out fe_tanh Vc=0.3498440821537202 Qo=1.2335190033420976e-13 K=2.62 tau=9.409402090143806e-08 off=-0.2

*Grain_748:
XU_748 in out fe_tanh Vc=0.18215990945546695 Qo=6.422795794546641e-14 K=2.62 tau=1.0733336881913872e-07 off=-0.2

*Grain_749:
XU_749 in out fe_tanh Vc=0.3563843701699473 Qo=1.2565794750404634e-13 K=2.62 tau=1.0469558354036783e-07 off=-0.2

*Grain_750:
XU_750 in out fe_tanh Vc=0.33383043851699634 Qo=1.1770563254055656e-13 K=2.62 tau=9.309544389242206e-08 off=-0.2

*Grain_751:
XU_751 in out fe_tanh Vc=0.24824988787743432 Qo=8.75306943565242e-14 K=2.62 tau=1.0954644784102406e-07 off=-0.2

*Grain_752:
XU_752 in out fe_tanh Vc=0.5885258361295903 Qo=2.0750895609109195e-13 K=2.62 tau=1.0095192640078747e-07 off=-0.2

*Grain_753:
XU_753 in out fe_tanh Vc=0.5649855534828199 Qo=1.9920886257226642e-13 K=2.62 tau=1.1082190475733947e-07 off=-0.2

*Grain_754:
XU_754 in out fe_tanh Vc=-0.22145767065991778 Qo=7.80839977378418e-14 K=2.62 tau=7.710770913029821e-08 off=-0.2

*Grain_755:
XU_755 in out fe_tanh Vc=0.9959127913304877 Qo=3.5114995978060915e-13 K=2.62 tau=1.0586775945233118e-07 off=-0.2

*Grain_756:
XU_756 in out fe_tanh Vc=0.48303691851057706 Qo=1.7031450543067847e-13 K=2.62 tau=9.117363768360323e-08 off=-0.2

*Grain_757:
XU_757 in out fe_tanh Vc=0.3254518761363255 Qo=1.1475142623996134e-13 K=2.62 tau=8.995140406682786e-08 off=-0.2

*Grain_758:
XU_758 in out fe_tanh Vc=0.6149455241630961 Qo=2.1682430224503365e-13 K=2.62 tau=9.57448417237228e-08 off=-0.2

*Grain_759:
XU_759 in out fe_tanh Vc=0.1012228810526824 Qo=3.5690284249729656e-14 K=2.62 tau=9.01648071639046e-08 off=-0.2

*Grain_760:
XU_760 in out fe_tanh Vc=0.6067372128681188 Qo=2.1393012495743466e-13 K=2.62 tau=9.106322204264256e-08 off=-0.2

*Grain_761:
XU_761 in out fe_tanh Vc=0.3644455594984296 Qo=1.2850025089960653e-13 K=2.62 tau=8.835294722784823e-08 off=-0.2

*Grain_762:
XU_762 in out fe_tanh Vc=0.7568314686881893 Qo=2.6685201967886534e-13 K=2.62 tau=9.508672829046297e-08 off=-0.2

*Grain_763:
XU_763 in out fe_tanh Vc=0.25453913905899067 Qo=8.974822817944384e-14 K=2.62 tau=9.661702807101889e-08 off=-0.2

*Grain_764:
XU_764 in out fe_tanh Vc=-0.0018849712944671304 Qo=6.646240514246849e-16 K=2.62 tau=9.485611303519025e-08 off=-0.2

*Grain_765:
XU_765 in out fe_tanh Vc=0.38716948127217016 Qo=1.3651250286219706e-13 K=2.62 tau=9.032230253959293e-08 off=-0.2

*Grain_766:
XU_766 in out fe_tanh Vc=0.7697073765328216 Qo=2.713919498425709e-13 K=2.62 tau=7.958355652063555e-08 off=-0.2

*Grain_767:
XU_767 in out fe_tanh Vc=0.6800147891397901 Qo=2.3976714420712423e-13 K=2.62 tau=9.243713708100012e-08 off=-0.2

*Grain_768:
XU_768 in out fe_tanh Vc=0.24341731728270077 Qo=8.58267731048345e-14 K=2.62 tau=9.896537265486608e-08 off=-0.2

*Grain_769:
XU_769 in out fe_tanh Vc=0.218218635010111 Qo=7.694194268236036e-14 K=2.62 tau=9.258248489177247e-08 off=-0.2

*Grain_770:
XU_770 in out fe_tanh Vc=0.5221255543249419 Qo=1.84096809477357e-13 K=2.62 tau=1.1700735798524423e-07 off=-0.2

*Grain_771:
XU_771 in out fe_tanh Vc=0.7017939571620235 Qo=2.4744628443068277e-13 K=2.62 tau=1.0437773053280732e-07 off=-0.2

*Grain_772:
XU_772 in out fe_tanh Vc=0.7898150976577714 Qo=2.784817528110345e-13 K=2.62 tau=9.823833551511754e-08 off=-0.2

*Grain_773:
XU_773 in out fe_tanh Vc=0.1740468588856563 Qo=6.136736873917548e-14 K=2.62 tau=9.683734734487023e-08 off=-0.2

*Grain_774:
XU_774 in out fe_tanh Vc=0.2102067025662413 Qo=7.411700682460191e-14 K=2.62 tau=1.0028332026452146e-07 off=-0.2

*Grain_775:
XU_775 in out fe_tanh Vc=0.46504691712561264 Qo=1.6397139153780045e-13 K=2.62 tau=1.0135282214302351e-07 off=-0.2

*Grain_776:
XU_776 in out fe_tanh Vc=0.9086999489210718 Qo=3.203994900898786e-13 K=2.62 tau=1.1303734816265036e-07 off=-0.2

*Grain_777:
XU_777 in out fe_tanh Vc=0.21406099706716933 Qo=7.547599665861678e-14 K=2.62 tau=1.0088539689987126e-07 off=-0.2

*Grain_778:
XU_778 in out fe_tanh Vc=0.27656451165887064 Qo=9.751417793922981e-14 K=2.62 tau=8.954493135609315e-08 off=-0.2

*Grain_779:
XU_779 in out fe_tanh Vc=0.8247911304956894 Qo=2.908139897611316e-13 K=2.62 tau=1.1216689234774417e-07 off=-0.2

*Grain_780:
XU_780 in out fe_tanh Vc=0.8995870653633917 Qo=3.1718636869750277e-13 K=2.62 tau=9.954657807038068e-08 off=-0.2

*Grain_781:
XU_781 in out fe_tanh Vc=0.4099970899368782 Qo=1.4456131389693722e-13 K=2.62 tau=1.1632304495219802e-07 off=-0.2

*Grain_782:
XU_782 in out fe_tanh Vc=0.45018920310642 Qo=1.5873269420838744e-13 K=2.62 tau=9.581114973625382e-08 off=-0.2

*Grain_783:
XU_783 in out fe_tanh Vc=1.3077566606185473 Qo=4.611033242835794e-13 K=2.62 tau=1.0467529931843835e-07 off=-0.2

*Grain_784:
XU_784 in out fe_tanh Vc=0.5703541245664532 Qo=2.0110177281150402e-13 K=2.62 tau=9.435771409093019e-08 off=-0.2

*Grain_785:
XU_785 in out fe_tanh Vc=0.3568773857712685 Qo=1.2583178040395705e-13 K=2.62 tau=1.1073824813579951e-07 off=-0.2

*Grain_786:
XU_786 in out fe_tanh Vc=0.7595676266234164 Qo=2.678167645413395e-13 K=2.62 tau=1.0520639289210961e-07 off=-0.2

*Grain_787:
XU_787 in out fe_tanh Vc=0.9366901272244139 Qo=3.3026857709330984e-13 K=2.62 tau=9.111973328103567e-08 off=-0.2

*Grain_788:
XU_788 in out fe_tanh Vc=-0.15153524598099338 Qo=5.342997498855559e-14 K=2.62 tau=1.0274840371234854e-07 off=-0.2

*Grain_789:
XU_789 in out fe_tanh Vc=-0.21378225969259862 Qo=7.537771634861182e-14 K=2.62 tau=8.792740005028526e-08 off=-0.2

*Grain_790:
XU_790 in out fe_tanh Vc=0.1302159551372788 Qo=4.5912983352852e-14 K=2.62 tau=1.1784318497422665e-07 off=-0.2

*Grain_791:
XU_791 in out fe_tanh Vc=0.3908379382628109 Qo=1.3780596804904283e-13 K=2.62 tau=8.876003551122127e-08 off=-0.2

*Grain_792:
XU_792 in out fe_tanh Vc=0.5671949801651375 Qo=1.9998788669705706e-13 K=2.62 tau=9.606968557359572e-08 off=-0.2

*Grain_793:
XU_793 in out fe_tanh Vc=0.21961501865564412 Qo=7.743429509035804e-14 K=2.62 tau=9.31011640902888e-08 off=-0.2

*Grain_794:
XU_794 in out fe_tanh Vc=0.5840578632613245 Qo=2.0593358874301683e-13 K=2.62 tau=8.537048516367804e-08 off=-0.2

*Grain_795:
XU_795 in out fe_tanh Vc=0.19270263490131467 Qo=6.794522882351351e-14 K=2.62 tau=9.293898212920467e-08 off=-0.2

*Grain_796:
XU_796 in out fe_tanh Vc=0.24147992889724665 Qo=8.514366725505142e-14 K=2.62 tau=1.1662622793569115e-07 off=-0.2

*Grain_797:
XU_797 in out fe_tanh Vc=1.0848241866326298 Qo=3.8249932405845425e-13 K=2.62 tau=9.962735226061179e-08 off=-0.2

*Grain_798:
XU_798 in out fe_tanh Vc=0.5993748089279566 Qo=2.113342070517888e-13 K=2.62 tau=8.937580013589073e-08 off=-0.2

*Grain_799:
XU_799 in out fe_tanh Vc=0.5641952613082508 Qo=1.9893021260639529e-13 K=2.62 tau=8.011302562605852e-08 off=-0.2

*Grain_800:
XU_800 in out fe_tanh Vc=0.7796754436740607 Qo=2.7490660133234673e-13 K=2.62 tau=9.52696930027831e-08 off=-0.2

*Grain_801:
XU_801 in out fe_tanh Vc=0.2083143719737351 Qo=7.344978795038458e-14 K=2.62 tau=1.1360401004926399e-07 off=-0.2

*Grain_802:
XU_802 in out fe_tanh Vc=0.7797236714691428 Qo=2.749236060223666e-13 K=2.62 tau=1.1169100993243018e-07 off=-0.2

*Grain_803:
XU_803 in out fe_tanh Vc=0.5205266665396157 Qo=1.835330559174083e-13 K=2.62 tau=8.451567989548588e-08 off=-0.2

*Grain_804:
XU_804 in out fe_tanh Vc=0.5115566854824085 Qo=1.8037032067101878e-13 K=2.62 tau=1.0500044107265998e-07 off=-0.2

*Grain_805:
XU_805 in out fe_tanh Vc=0.5239913142625809 Qo=1.8475465977586252e-13 K=2.62 tau=1.0025693268815592e-07 off=-0.2

*Grain_806:
XU_806 in out fe_tanh Vc=0.5425509899946729 Qo=1.912986357580954e-13 K=2.62 tau=1.1625238628900368e-07 off=-0.2

*Grain_807:
XU_807 in out fe_tanh Vc=0.18005996865325896 Qo=6.348753756462977e-14 K=2.62 tau=9.811790837534565e-08 off=-0.2

*Grain_808:
XU_808 in out fe_tanh Vc=0.7917970073199029 Qo=2.7918055646553573e-13 K=2.62 tau=1.0174713111986571e-07 off=-0.2

*Grain_809:
XU_809 in out fe_tanh Vc=0.16808761938227734 Qo=5.926619408799045e-14 K=2.62 tau=1.1782189150629147e-07 off=-0.2

*Grain_810:
XU_810 in out fe_tanh Vc=0.2503959130321053 Qo=8.828736366864755e-14 K=2.62 tau=1.0323744045581484e-07 off=-0.2

*Grain_811:
XU_811 in out fe_tanh Vc=0.07403353956565095 Qo=2.6103565158716352e-14 K=2.62 tau=1.1076561407111805e-07 off=-0.2

*Grain_812:
XU_812 in out fe_tanh Vc=0.3815817022694286 Qo=1.3454230186753536e-13 K=2.62 tau=1.0560556643569419e-07 off=-0.2

*Grain_813:
XU_813 in out fe_tanh Vc=1.4704755556765483 Qo=5.184765541010495e-13 K=2.62 tau=1.0130963078649149e-07 off=-0.2

*Grain_814:
XU_814 in out fe_tanh Vc=0.17703313675372612 Qo=6.242030365716716e-14 K=2.62 tau=1.0394728562776817e-07 off=-0.2

*Grain_815:
XU_815 in out fe_tanh Vc=0.8315691596204523 Qo=2.9320386232354e-13 K=2.62 tau=1.0306715386562027e-07 off=-0.2

*Grain_816:
XU_816 in out fe_tanh Vc=0.8522154091748362 Qo=3.004835456088172e-13 K=2.62 tau=9.705340665523063e-08 off=-0.2

*Grain_817:
XU_817 in out fe_tanh Vc=0.5300168563704476 Qo=1.8687921213351129e-13 K=2.62 tau=9.395955681821256e-08 off=-0.2

*Grain_818:
XU_818 in out fe_tanh Vc=0.722705973930478 Qo=2.5481967486315627e-13 K=2.62 tau=9.218145204891199e-08 off=-0.2

*Grain_819:
XU_819 in out fe_tanh Vc=0.22314780384569521 Qo=7.86799236114484e-14 K=2.62 tau=9.110363046787334e-08 off=-0.2

*Grain_820:
XU_820 in out fe_tanh Vc=0.3203724725129277 Qo=1.1296047386582548e-13 K=2.62 tau=9.805714499616856e-08 off=-0.2

*Grain_821:
XU_821 in out fe_tanh Vc=0.7257467360736065 Qo=2.5589182045015643e-13 K=2.62 tau=1.112612073477072e-07 off=-0.2

*Grain_822:
XU_822 in out fe_tanh Vc=0.2801991627569838 Qo=9.879572347015316e-14 K=2.62 tau=9.237128456258189e-08 off=-0.2

*Grain_823:
XU_823 in out fe_tanh Vc=0.22997303914405215 Qo=8.108644064925991e-14 K=2.62 tau=1.1351439321345692e-07 off=-0.2

*Grain_824:
XU_824 in out fe_tanh Vc=1.1109111835431087 Qo=3.9169736629232663e-13 K=2.62 tau=1.2720390235140548e-07 off=-0.2

*Grain_825:
XU_825 in out fe_tanh Vc=1.392813686151045 Qo=4.910936721883321e-13 K=2.62 tau=1.0153548791609555e-07 off=-0.2

*Grain_826:
XU_826 in out fe_tanh Vc=0.5465244682475764 Qo=1.9269964871911196e-13 K=2.62 tau=9.617695286088415e-08 off=-0.2

*Grain_827:
XU_827 in out fe_tanh Vc=0.2963840392995546 Qo=1.0450236645782403e-13 K=2.62 tau=1.3119919709918354e-07 off=-0.2

*Grain_828:
XU_828 in out fe_tanh Vc=0.5250569216683819 Qo=1.8513038343454657e-13 K=2.62 tau=8.680732414840708e-08 off=-0.2

*Grain_829:
XU_829 in out fe_tanh Vc=0.576330349766193 Qo=2.032089364675958e-13 K=2.62 tau=1.0052709169938832e-07 off=-0.2

*Grain_830:
XU_830 in out fe_tanh Vc=1.3893144035142837 Qo=4.898598563684569e-13 K=2.62 tau=1.0503209302981141e-07 off=-0.2

*Grain_831:
XU_831 in out fe_tanh Vc=0.829305106166681 Qo=2.924055772867841e-13 K=2.62 tau=1.0488717405970469e-07 off=-0.2

*Grain_832:
XU_832 in out fe_tanh Vc=0.606276463012335 Qo=2.1376766867136642e-13 K=2.62 tau=8.564463753725216e-08 off=-0.2

*Grain_833:
XU_833 in out fe_tanh Vc=0.38301621778928885 Qo=1.3504809923402026e-13 K=2.62 tau=1.0629520223542859e-07 off=-0.2

*Grain_834:
XU_834 in out fe_tanh Vc=0.09713176919302624 Qo=3.4247794729078936e-14 K=2.62 tau=9.639089560298312e-08 off=-0.2

*Grain_835:
XU_835 in out fe_tanh Vc=0.602246229435176 Qo=2.1234664428966813e-13 K=2.62 tau=1.1053112173731112e-07 off=-0.2

*Grain_836:
XU_836 in out fe_tanh Vc=0.8436728821332777 Qo=2.974715268324939e-13 K=2.62 tau=1.0729385717477861e-07 off=-0.2

*Grain_837:
XU_837 in out fe_tanh Vc=0.26214275665183473 Qo=9.242919586572822e-14 K=2.62 tau=1.1137001973156448e-07 off=-0.2

*Grain_838:
XU_838 in out fe_tanh Vc=0.6560864139587972 Qo=2.313302127252063e-13 K=2.62 tau=1.140311936481691e-07 off=-0.2

*Grain_839:
XU_839 in out fe_tanh Vc=-0.0763461833054338 Qo=2.6918982696557913e-14 K=2.62 tau=9.557899034337256e-08 off=-0.2

*Grain_840:
XU_840 in out fe_tanh Vc=0.5031199569033818 Qo=1.773956054881288e-13 K=2.62 tau=1.2247507600243363e-07 off=-0.2

*Grain_841:
XU_841 in out fe_tanh Vc=1.0066497704857813 Qo=3.549357227825178e-13 K=2.62 tau=1.142817914593603e-07 off=-0.2

*Grain_842:
XU_842 in out fe_tanh Vc=0.8086046949761638 Qo=2.8510679709210336e-13 K=2.62 tau=1.092953294740162e-07 off=-0.2

*Grain_843:
XU_843 in out fe_tanh Vc=0.2119483207244493 Qo=7.473108583988486e-14 K=2.62 tau=9.193240652161875e-08 off=-0.2

*Grain_844:
XU_844 in out fe_tanh Vc=0.7940822318367391 Qo=2.799863062301358e-13 K=2.62 tau=1.0997130585071424e-07 off=-0.2

*Grain_845:
XU_845 in out fe_tanh Vc=0.5046789229622428 Qo=1.7794528300370425e-13 K=2.62 tau=1.0263721954379955e-07 off=-0.2

*Grain_846:
XU_846 in out fe_tanh Vc=0.6545766554374018 Qo=2.30797885348069e-13 K=2.62 tau=1.1367223474800125e-07 off=-0.2

*Grain_847:
XU_847 in out fe_tanh Vc=0.9660821683945136 Qo=3.406319484292299e-13 K=2.62 tau=1.0546336325413309e-07 off=-0.2

*Grain_848:
XU_848 in out fe_tanh Vc=0.20471943891326766 Qo=7.218224664497502e-14 K=2.62 tau=8.514265791178012e-08 off=-0.2

*Grain_849:
XU_849 in out fe_tanh Vc=0.4625324040766766 Qo=1.630847966836244e-13 K=2.62 tau=1.1385551175185018e-07 off=-0.2

*Grain_850:
XU_850 in out fe_tanh Vc=0.5016985383318892 Qo=1.7689442598872276e-13 K=2.62 tau=9.369544107962121e-08 off=-0.2

*Grain_851:
XU_851 in out fe_tanh Vc=0.5091128381958494 Qo=1.7950864193382862e-13 K=2.62 tau=9.324706613255941e-08 off=-0.2

*Grain_852:
XU_852 in out fe_tanh Vc=0.02567388219981015 Qo=9.052381674736146e-15 K=2.62 tau=1.2242426093803727e-07 off=-0.2

*Grain_853:
XU_853 in out fe_tanh Vc=0.3829389973096332 Qo=1.3502087198223537e-13 K=2.62 tau=1.1168170294446949e-07 off=-0.2

*Grain_854:
XU_854 in out fe_tanh Vc=0.2495621862259698 Qo=8.799339903942396e-14 K=2.62 tau=9.388904652489026e-08 off=-0.2

*Grain_855:
XU_855 in out fe_tanh Vc=0.6112274521691621 Qo=2.1551334325093627e-13 K=2.62 tau=9.480292369230388e-08 off=-0.2

*Grain_856:
XU_856 in out fe_tanh Vc=0.23386103601333086 Qo=8.245731363749659e-14 K=2.62 tau=9.66489822428673e-08 off=-0.2

*Grain_857:
XU_857 in out fe_tanh Vc=1.2185220103619685 Qo=4.2963998319447374e-13 K=2.62 tau=1.105229492245877e-07 off=-0.2

*Grain_858:
XU_858 in out fe_tanh Vc=0.4291102141106447 Qo=1.5130043085910977e-13 K=2.62 tau=1.2019276656487896e-07 off=-0.2

*Grain_859:
XU_859 in out fe_tanh Vc=0.4468459415459614 Qo=1.5755389002722743e-13 K=2.62 tau=9.12985051421697e-08 off=-0.2

*Grain_860:
XU_860 in out fe_tanh Vc=0.1751856713136189 Qo=6.176890383517769e-14 K=2.62 tau=1.0813519118355846e-07 off=-0.2

*Grain_861:
XU_861 in out fe_tanh Vc=0.19573390067073887 Qo=6.901402607391896e-14 K=2.62 tau=1.0722741099218279e-07 off=-0.2

*Grain_862:
XU_862 in out fe_tanh Vc=0.7475459574120287 Qo=2.6357803129398855e-13 K=2.62 tau=9.318144556981908e-08 off=-0.2

*Grain_863:
XU_863 in out fe_tanh Vc=0.15090775881589247 Qo=5.3208728615674215e-14 K=2.62 tau=1.14804577149126e-07 off=-0.2

*Grain_864:
XU_864 in out fe_tanh Vc=1.0029688454319625 Qo=3.5363786146789703e-13 K=2.62 tau=1.1703511427188191e-07 off=-0.2

*Grain_865:
XU_865 in out fe_tanh Vc=0.35753596577070496 Qo=1.2606398983266165e-13 K=2.62 tau=1.0142290948514324e-07 off=-0.2

*Grain_866:
XU_866 in out fe_tanh Vc=0.8140092401379848 Qo=2.8701239147017186e-13 K=2.62 tau=9.657306202298633e-08 off=-0.2

*Grain_867:
XU_867 in out fe_tanh Vc=0.06978320326067589 Qo=2.4604934520031465e-14 K=2.62 tau=1.0771103116877614e-07 off=-0.2

*Grain_868:
XU_868 in out fe_tanh Vc=0.8142938169314926 Qo=2.87112730707166e-13 K=2.62 tau=8.659297681276843e-08 off=-0.2

*Grain_869:
XU_869 in out fe_tanh Vc=0.15424631496061886 Qo=5.4385873709251935e-14 K=2.62 tau=7.701336980757947e-08 off=-0.2

*Grain_870:
XU_870 in out fe_tanh Vc=0.498837960691757 Qo=1.7588581184898493e-13 K=2.62 tau=8.432385293743638e-08 off=-0.2

*Grain_871:
XU_871 in out fe_tanh Vc=0.6052278070174959 Qo=2.133979219288635e-13 K=2.62 tau=9.787516036647695e-08 off=-0.2

*Grain_872:
XU_872 in out fe_tanh Vc=0.8743456103579088 Qo=3.082864569912396e-13 K=2.62 tau=1.0093725016363249e-07 off=-0.2

*Grain_873:
XU_873 in out fe_tanh Vc=0.1924227724719395 Qo=6.784655182922779e-14 K=2.62 tau=1.0473084202218354e-07 off=-0.2

*Grain_874:
XU_874 in out fe_tanh Vc=0.7756543758419628 Qo=2.73488808710535e-13 K=2.62 tau=1.0112057653000082e-07 off=-0.2

*Grain_875:
XU_875 in out fe_tanh Vc=0.5224361379553488 Qo=1.8420631849288054e-13 K=2.62 tau=1.0029371494963031e-07 off=-0.2

*Grain_876:
XU_876 in out fe_tanh Vc=0.48474727097599374 Qo=1.709175604417898e-13 K=2.62 tau=9.991025466820008e-08 off=-0.2

*Grain_877:
XU_877 in out fe_tanh Vc=0.5204302101850183 Qo=1.8349904626783628e-13 K=2.62 tau=1.1647017734889801e-07 off=-0.2

*Grain_878:
XU_878 in out fe_tanh Vc=0.4392972509320286 Qo=1.548922891033779e-13 K=2.62 tau=1.1248016593059661e-07 off=-0.2

*Grain_879:
XU_879 in out fe_tanh Vc=0.9886035717581934 Qo=3.4857279420830036e-13 K=2.62 tau=1.0446967100643641e-07 off=-0.2

*Grain_880:
XU_880 in out fe_tanh Vc=0.021804722767279017 Qo=7.688150598536212e-15 K=2.62 tau=1.03380732625476e-07 off=-0.2

*Grain_881:
XU_881 in out fe_tanh Vc=0.3489085181044919 Qo=1.2302202880216547e-13 K=2.62 tau=1.0380343332807141e-07 off=-0.2

*Grain_882:
XU_882 in out fe_tanh Vc=0.19475138916549212 Qo=6.866760128797915e-14 K=2.62 tau=1.0675383109555271e-07 off=-0.2

*Grain_883:
XU_883 in out fe_tanh Vc=0.6578569387005018 Qo=2.3195448394378313e-13 K=2.62 tau=1.1129556666459872e-07 off=-0.2

*Grain_884:
XU_884 in out fe_tanh Vc=0.45490090824103 Qo=1.6039399937779493e-13 K=2.62 tau=9.783822843783624e-08 off=-0.2

*Grain_885:
XU_885 in out fe_tanh Vc=0.2979613807339976 Qo=1.0505852296679405e-13 K=2.62 tau=1.0917328046059888e-07 off=-0.2

*Grain_886:
XU_886 in out fe_tanh Vc=0.09058711861547919 Qo=3.1940209359065194e-14 K=2.62 tau=1.0796141685961772e-07 off=-0.2

*Grain_887:
XU_887 in out fe_tanh Vc=0.9753612267847225 Qo=3.4390366158412453e-13 K=2.62 tau=8.967133896804752e-08 off=-0.2

*Grain_888:
XU_888 in out fe_tanh Vc=0.46009114484353403 Qo=1.6222403047096554e-13 K=2.62 tau=1.0806946005295761e-07 off=-0.2

*Grain_889:
XU_889 in out fe_tanh Vc=0.5196990434051526 Qo=1.8324124338832938e-13 K=2.62 tau=1.0587743858451069e-07 off=-0.2

*Grain_890:
XU_890 in out fe_tanh Vc=0.7850928086684326 Qo=2.7681671586893094e-13 K=2.62 tau=9.968300610956435e-08 off=-0.2

*Grain_891:
XU_891 in out fe_tanh Vc=0.4283566815531913 Qo=1.5103474200608315e-13 K=2.62 tau=1.044192099410491e-07 off=-0.2

*Grain_892:
XU_892 in out fe_tanh Vc=0.2802951461511836 Qo=9.882956635811109e-14 K=2.62 tau=8.38186182012157e-08 off=-0.2

*Grain_893:
XU_893 in out fe_tanh Vc=0.24722087380949373 Qo=8.716787318210361e-14 K=2.62 tau=7.461874456640157e-08 off=-0.2

*Grain_894:
XU_894 in out fe_tanh Vc=-0.4005670343725572 Qo=1.4123636048639168e-13 K=2.62 tau=9.625870696319301e-08 off=-0.2

*Grain_895:
XU_895 in out fe_tanh Vc=0.09148809826757909 Qo=3.225788674141447e-14 K=2.62 tau=9.014200912693936e-08 off=-0.2

*Grain_896:
XU_896 in out fe_tanh Vc=0.4388027187839 Qo=1.54717921482601e-13 K=2.62 tau=9.381915856726934e-08 off=-0.2

*Grain_897:
XU_897 in out fe_tanh Vc=0.49051886883542883 Qo=1.729525743243838e-13 K=2.62 tau=9.518915622453776e-08 off=-0.2

*Grain_898:
XU_898 in out fe_tanh Vc=0.4207214359527056 Qo=1.4834262256664527e-13 K=2.62 tau=9.695860916808253e-08 off=-0.2

*Grain_899:
XU_899 in out fe_tanh Vc=0.40906852511036984 Qo=1.442339102283424e-13 K=2.62 tau=1.18538839424134e-07 off=-0.2

*Grain_900:
XU_900 in out fe_tanh Vc=0.5342367195448107 Qo=1.8836709821837383e-13 K=2.62 tau=9.317705692308071e-08 off=-0.2

*Grain_901:
XU_901 in out fe_tanh Vc=0.09351952216185433 Qo=3.2974148672159563e-14 K=2.62 tau=1.0223362378622606e-07 off=-0.2

*Grain_902:
XU_902 in out fe_tanh Vc=0.6768289694685813 Qo=2.3864385263064123e-13 K=2.62 tau=1.1417786983589754e-07 off=-0.2

*Grain_903:
XU_903 in out fe_tanh Vc=0.6161985386819182 Qo=2.17266103978799e-13 K=2.62 tau=9.152754759469263e-08 off=-0.2

*Grain_904:
XU_904 in out fe_tanh Vc=0.3722268090036822 Qo=1.3124385001249874e-13 K=2.62 tau=1.1421225009284181e-07 off=-0.2

*Grain_905:
XU_905 in out fe_tanh Vc=0.41107864572562847 Qo=1.449426608130791e-13 K=2.62 tau=9.690603956838706e-08 off=-0.2

*Grain_906:
XU_906 in out fe_tanh Vc=0.5456964034822331 Qo=1.924076804749271e-13 K=2.62 tau=9.550739931203642e-08 off=-0.2

*Grain_907:
XU_907 in out fe_tanh Vc=0.11810774781013927 Qo=4.16437375384066e-14 K=2.62 tau=1.0632873153556516e-07 off=-0.2

*Grain_908:
XU_908 in out fe_tanh Vc=0.7386869188335459 Qo=2.6045441337522165e-13 K=2.62 tau=1.2469965465489444e-07 off=-0.2

*Grain_909:
XU_909 in out fe_tanh Vc=0.8141792194243644 Qo=2.870723246491564e-13 K=2.62 tau=9.627818879812825e-08 off=-0.2

*Grain_910:
XU_910 in out fe_tanh Vc=0.42431196547084193 Qo=1.4960861122233898e-13 K=2.62 tau=1.2405064246831793e-07 off=-0.2

*Grain_911:
XU_911 in out fe_tanh Vc=0.3295700302393805 Qo=1.1620345061423032e-13 K=2.62 tau=8.794353255366338e-08 off=-0.2

*Grain_912:
XU_912 in out fe_tanh Vc=0.49808800570352096 Qo=1.7562138441492765e-13 K=2.62 tau=9.553429905161607e-08 off=-0.2

*Grain_913:
XU_913 in out fe_tanh Vc=0.26291993437749434 Qo=9.270322179398562e-14 K=2.62 tau=1.0022712404154226e-07 off=-0.2

*Grain_914:
XU_914 in out fe_tanh Vc=0.48617014429384586 Qo=1.7141925287177574e-13 K=2.62 tau=1.0372625150328708e-07 off=-0.2

*Grain_915:
XU_915 in out fe_tanh Vc=0.3542983756760943 Qo=1.24922444467038e-13 K=2.62 tau=7.870645542456462e-08 off=-0.2

*Grain_916:
XU_916 in out fe_tanh Vc=0.6916609654687115 Qo=2.4387348201611575e-13 K=2.62 tau=9.361763438238374e-08 off=-0.2

*Grain_917:
XU_917 in out fe_tanh Vc=0.4932967914593822 Qo=1.7393204504327247e-13 K=2.62 tau=8.877168883686634e-08 off=-0.2

*Grain_918:
XU_918 in out fe_tanh Vc=0.07030284821308597 Qo=2.4788156691417797e-14 K=2.62 tau=9.007039242988153e-08 off=-0.2

*Grain_919:
XU_919 in out fe_tanh Vc=0.5616183991735114 Qo=1.9802163402115086e-13 K=2.62 tau=1.0412395166245334e-07 off=-0.2

*Grain_920:
XU_920 in out fe_tanh Vc=0.8032286195604593 Qo=2.8321124089236813e-13 K=2.62 tau=9.518860943554498e-08 off=-0.2

*Grain_921:
XU_921 in out fe_tanh Vc=0.402509673790978 Qo=1.419213178035232e-13 K=2.62 tau=9.901476082120366e-08 off=-0.2

*Grain_922:
XU_922 in out fe_tanh Vc=0.874679701218094 Qo=3.0840425444613564e-13 K=2.62 tau=8.157256395946343e-08 off=-0.2

*Grain_923:
XU_923 in out fe_tanh Vc=0.6361015526066074 Qo=2.2428372901585735e-13 K=2.62 tau=1.016317547796172e-07 off=-0.2

*Grain_924:
XU_924 in out fe_tanh Vc=0.42799122240655274 Qo=1.5090588437340613e-13 K=2.62 tau=9.760183584128143e-08 off=-0.2

*Grain_925:
XU_925 in out fe_tanh Vc=0.19268020799634594 Qo=6.793732129702493e-14 K=2.62 tau=9.221867924617849e-08 off=-0.2

*Grain_926:
XU_926 in out fe_tanh Vc=0.2830201415740159 Qo=9.979037541836179e-14 K=2.62 tau=1.1673051851564253e-07 off=-0.2

*Grain_927:
XU_927 in out fe_tanh Vc=-0.19986604567372895 Qo=7.047098351460928e-14 K=2.62 tau=1.0565663252100603e-07 off=-0.2

*Grain_928:
XU_928 in out fe_tanh Vc=0.19617496780046578 Qo=6.916954240648583e-14 K=2.62 tau=1.0646506544017842e-07 off=-0.2

*Grain_929:
XU_929 in out fe_tanh Vc=0.5388507494362325 Qo=1.8999396396897313e-13 K=2.62 tau=1.0464033661046777e-07 off=-0.2

*Grain_930:
XU_930 in out fe_tanh Vc=0.3437574382463031 Qo=1.2120580402749093e-13 K=2.62 tau=9.443599191584848e-08 off=-0.2

*Grain_931:
XU_931 in out fe_tanh Vc=-0.1717222234692512 Qo=6.054772304320575e-14 K=2.62 tau=1.093598349284638e-07 off=-0.2

*Grain_932:
XU_932 in out fe_tanh Vc=1.0879212691671845 Qo=3.8359132771270317e-13 K=2.62 tau=1.0418291214508417e-07 off=-0.2

*Grain_933:
XU_933 in out fe_tanh Vc=0.14212314020494404 Qo=5.011135051311816e-14 K=2.62 tau=8.342459774536728e-08 off=-0.2

*Grain_934:
XU_934 in out fe_tanh Vc=0.22006396790282257 Qo=7.759259058717522e-14 K=2.62 tau=1.1460377598343612e-07 off=-0.2

*Grain_935:
XU_935 in out fe_tanh Vc=0.3518389882157271 Qo=1.2405528640328915e-13 K=2.62 tau=9.921201300425912e-08 off=-0.2

*Grain_936:
XU_936 in out fe_tanh Vc=0.46258888681658056 Qo=1.6310471199349715e-13 K=2.62 tau=1.0146174690443866e-07 off=-0.2

*Grain_937:
XU_937 in out fe_tanh Vc=0.8233302253714117 Qo=2.9029888765570726e-13 K=2.62 tau=9.719656870783383e-08 off=-0.2

*Grain_938:
XU_938 in out fe_tanh Vc=-0.07103782503803063 Qo=2.5047302958807543e-14 K=2.62 tau=1.1438240885226278e-07 off=-0.2

*Grain_939:
XU_939 in out fe_tanh Vc=1.2750754783435752 Qo=4.4958023115600955e-13 K=2.62 tau=9.330593461279377e-08 off=-0.2

*Grain_940:
XU_940 in out fe_tanh Vc=0.2841693561336613 Qo=1.0019557821313628e-13 K=2.62 tau=1.0339209649104597e-07 off=-0.2

*Grain_941:
XU_941 in out fe_tanh Vc=0.16644902918691434 Qo=5.868844181268338e-14 K=2.62 tau=9.274534464370725e-08 off=-0.2

*Grain_942:
XU_942 in out fe_tanh Vc=0.9112807666794197 Qo=3.2130946339269587e-13 K=2.62 tau=1.1173147174713515e-07 off=-0.2

*Grain_943:
XU_943 in out fe_tanh Vc=0.7645970238318869 Qo=2.695900850999757e-13 K=2.62 tau=1.0854302741612962e-07 off=-0.2

*Grain_944:
XU_944 in out fe_tanh Vc=0.39863908365020834 Qo=1.4055658227237017e-13 K=2.62 tau=1.0918395338590765e-07 off=-0.2

*Grain_945:
XU_945 in out fe_tanh Vc=0.05238159043720486 Qo=1.846928118143324e-14 K=2.62 tau=9.344321584910501e-08 off=-0.2

*Grain_946:
XU_946 in out fe_tanh Vc=0.6126269810269789 Qo=2.1600680463270807e-13 K=2.62 tau=1.0536672046100535e-07 off=-0.2

*Grain_947:
XU_947 in out fe_tanh Vc=0.7570834819149035 Qo=2.6694087729290066e-13 K=2.62 tau=9.785406873468621e-08 off=-0.2

*Grain_948:
XU_948 in out fe_tanh Vc=0.30648635186829437 Qo=1.0806435168693726e-13 K=2.62 tau=9.997094382912027e-08 off=-0.2

*Grain_949:
XU_949 in out fe_tanh Vc=0.43925538445428514 Qo=1.5487752735706464e-13 K=2.62 tau=9.6149905522889e-08 off=-0.2

*Grain_950:
XU_950 in out fe_tanh Vc=0.39439054823759456 Qo=1.3905858661225545e-13 K=2.62 tau=8.984909439718147e-08 off=-0.2

*Grain_951:
XU_951 in out fe_tanh Vc=0.2068238663563283 Qo=7.292424897532437e-14 K=2.62 tau=7.315404462045866e-08 off=-0.2

*Grain_952:
XU_952 in out fe_tanh Vc=0.466372692572275 Qo=1.6443884812519064e-13 K=2.62 tau=1.0894254017640606e-07 off=-0.2

*Grain_953:
XU_953 in out fe_tanh Vc=1.1222732751533802 Qo=3.9570353836552616e-13 K=2.62 tau=8.852894268446706e-08 off=-0.2

*Grain_954:
XU_954 in out fe_tanh Vc=0.6617141391807473 Qo=2.3331449840016385e-13 K=2.62 tau=1.0893709095294133e-07 off=-0.2

*Grain_955:
XU_955 in out fe_tanh Vc=0.7163111369042441 Qo=2.525649124139607e-13 K=2.62 tau=7.893763414130185e-08 off=-0.2

*Grain_956:
XU_956 in out fe_tanh Vc=0.5386837896697959 Qo=1.899350954457655e-13 K=2.62 tau=9.875378317633131e-08 off=-0.2

*Grain_957:
XU_957 in out fe_tanh Vc=0.6862555814223422 Qo=2.4196759185484415e-13 K=2.62 tau=9.914343529655393e-08 off=-0.2

*Grain_958:
XU_958 in out fe_tanh Vc=-0.16086018139009434 Qo=5.671786397077067e-14 K=2.62 tau=1.0859934003659158e-07 off=-0.2

*Grain_959:
XU_959 in out fe_tanh Vc=0.9665646664830354 Qo=3.408020729480167e-13 K=2.62 tau=1.11319103288376e-07 off=-0.2

*Grain_960:
XU_960 in out fe_tanh Vc=0.10871206538731815 Qo=3.833090379070733e-14 K=2.62 tau=1.1221844204212398e-07 off=-0.2

*Grain_961:
XU_961 in out fe_tanh Vc=0.16861529760323501 Qo=5.945224871815426e-14 K=2.62 tau=8.466479436888942e-08 off=-0.2

*Grain_962:
XU_962 in out fe_tanh Vc=0.7796032390337323 Qo=2.748811426207326e-13 K=2.62 tau=8.53454957546178e-08 off=-0.2

*Grain_963:
XU_963 in out fe_tanh Vc=0.011124973204846511 Qo=3.9225662401858304e-15 K=2.62 tau=1.028752426386755e-07 off=-0.2

*Grain_964:
XU_964 in out fe_tanh Vc=1.1320507936190418 Qo=3.9915100409330785e-13 K=2.62 tau=9.568246907799934e-08 off=-0.2

*Grain_965:
XU_965 in out fe_tanh Vc=0.7052922741648104 Qo=2.486797597766388e-13 K=2.62 tau=1.0365840989753072e-07 off=-0.2

*Grain_966:
XU_966 in out fe_tanh Vc=0.631785182935978 Qo=2.227618156019179e-13 K=2.62 tau=1.0878232373923691e-07 off=-0.2

*Grain_967:
XU_967 in out fe_tanh Vc=0.5968394944389126 Qo=2.1044027779552367e-13 K=2.62 tau=9.649821446101897e-08 off=-0.2

*Grain_968:
XU_968 in out fe_tanh Vc=0.2703626431503139 Qo=9.532745446675095e-14 K=2.62 tau=1.0895480880138833e-07 off=-0.2

*Grain_969:
XU_969 in out fe_tanh Vc=0.8934793418992832 Qo=3.150328399272702e-13 K=2.62 tau=1.0201931356951208e-07 off=-0.2

*Grain_970:
XU_970 in out fe_tanh Vc=-0.129204843208035 Qo=4.555647431272478e-14 K=2.62 tau=9.321274170646448e-08 off=-0.2

*Grain_971:
XU_971 in out fe_tanh Vc=0.45361689291044494 Qo=1.5994126703454398e-13 K=2.62 tau=1.1822836747413925e-07 off=-0.2

*Grain_972:
XU_972 in out fe_tanh Vc=-0.586086840890043 Qo=2.066489881423643e-13 K=2.62 tau=9.325004017251217e-08 off=-0.2

*Grain_973:
XU_973 in out fe_tanh Vc=0.3298404862694515 Qo=1.1629881099609165e-13 K=2.62 tau=9.322984712988239e-08 off=-0.2

*Grain_974:
XU_974 in out fe_tanh Vc=0.28431254303331044 Qo=1.0024606463573331e-13 K=2.62 tau=1.0437066326655952e-07 off=-0.2

*Grain_975:
XU_975 in out fe_tanh Vc=0.020177785212107557 Qo=7.114506940138378e-15 K=2.62 tau=1.0569524996718025e-07 off=-0.2

*Grain_976:
XU_976 in out fe_tanh Vc=0.29709260482405186 Qo=1.0475220033644783e-13 K=2.62 tau=1.1033941893500247e-07 off=-0.2

*Grain_977:
XU_977 in out fe_tanh Vc=0.7230782298528676 Qo=2.549509289782888e-13 K=2.62 tau=1.0178768408484447e-07 off=-0.2

*Grain_978:
XU_978 in out fe_tanh Vc=1.2198790008792086 Qo=4.3011844593709497e-13 K=2.62 tau=9.512137165135107e-08 off=-0.2

*Grain_979:
XU_979 in out fe_tanh Vc=0.3747642652316991 Qo=1.3213853442680655e-13 K=2.62 tau=9.217734304879738e-08 off=-0.2

*Grain_980:
XU_980 in out fe_tanh Vc=0.4866616611048246 Qo=1.715925573115913e-13 K=2.62 tau=1.0272749380172013e-07 off=-0.2

*Grain_981:
XU_981 in out fe_tanh Vc=0.04233299670570595 Qo=1.4926236734786915e-14 K=2.62 tau=1.0326232807461744e-07 off=-0.2

*Grain_982:
XU_982 in out fe_tanh Vc=0.07105395640469364 Qo=2.505299073468936e-14 K=2.62 tau=1.048053008878689e-07 off=-0.2

*Grain_983:
XU_983 in out fe_tanh Vc=0.2427955640125066 Qo=8.560754845211117e-14 K=2.62 tau=8.226977602970326e-08 off=-0.2

*Grain_984:
XU_984 in out fe_tanh Vc=0.32327826855336333 Qo=1.139850316098489e-13 K=2.62 tau=9.312145850054283e-08 off=-0.2

*Grain_985:
XU_985 in out fe_tanh Vc=0.4082382083221307 Qo=1.439411479409881e-13 K=2.62 tau=1.0718637375843548e-07 off=-0.2

*Grain_986:
XU_986 in out fe_tanh Vc=0.5317784026781788 Qo=1.8750031763641892e-13 K=2.62 tau=1.0087607021146713e-07 off=-0.2

*Grain_987:
XU_987 in out fe_tanh Vc=0.5679502997346575 Qo=2.0025420563458584e-13 K=2.62 tau=9.76465933334587e-08 off=-0.2

*Grain_988:
XU_988 in out fe_tanh Vc=0.7845509804674076 Qo=2.766256720821113e-13 K=2.62 tau=7.224389759946893e-08 off=-0.2

*Grain_989:
XU_989 in out fe_tanh Vc=0.673093562619502 Qo=2.373267815213666e-13 K=2.62 tau=1.1317245693714194e-07 off=-0.2

*Grain_990:
XU_990 in out fe_tanh Vc=0.5165781419242768 Qo=1.8214084138623767e-13 K=2.62 tau=1.2184113625959763e-07 off=-0.2

*Grain_991:
XU_991 in out fe_tanh Vc=0.3332274911264356 Qo=1.1749303867311323e-13 K=2.62 tau=1.1655982296100885e-07 off=-0.2

*Grain_992:
XU_992 in out fe_tanh Vc=0.653950854536799 Qo=2.3057723353699655e-13 K=2.62 tau=9.958246285581624e-08 off=-0.2

*Grain_993:
XU_993 in out fe_tanh Vc=0.11277146251155074 Qo=3.9762210978762885e-14 K=2.62 tau=1.0329673873093171e-07 off=-0.2

*Grain_994:
XU_994 in out fe_tanh Vc=0.056601458836247676 Qo=1.995716910847124e-14 K=2.62 tau=1.2521091786060875e-07 off=-0.2

*Grain_995:
XU_995 in out fe_tanh Vc=0.32924123049830395 Qo=1.160875187606986e-13 K=2.62 tau=8.533277185756104e-08 off=-0.2

*Grain_996:
XU_996 in out fe_tanh Vc=0.15705559645831968 Qo=5.5376401287085496e-14 K=2.62 tau=1.0087280289994053e-07 off=-0.2

*Grain_997:
XU_997 in out fe_tanh Vc=0.5001048562601971 Qo=1.7633250791693044e-13 K=2.62 tau=9.681275717190352e-08 off=-0.2

*Grain_998:
XU_998 in out fe_tanh Vc=0.3738721400385161 Qo=1.3182397904762825e-13 K=2.62 tau=1.1110580688762471e-07 off=-0.2

*Grain_999:
XU_999 in out fe_tanh Vc=0.5400328272721624 Qo=1.9041075406159739e-13 K=2.62 tau=9.550669296252931e-08 off=-0.2

*Grain_1000:
XU_1000 in out fe_tanh Vc=0.5175852107807777 Qo=1.8249592487500796e-13 K=2.62 tau=9.843926446614918e-08 off=-0.2

*Grain_1001:
XU_1001 in out fe_tanh Vc=0.15975391512755172 Qo=5.632780436215823e-14 K=2.62 tau=1.1659359225850965e-07 off=-0.2

*Grain_1002:
XU_1002 in out fe_tanh Vc=-0.07136768238860819 Qo=2.5163607716008125e-14 K=2.62 tau=1.0600939092020414e-07 off=-0.2

*Grain_1003:
XU_1003 in out fe_tanh Vc=0.5579695006029444 Qo=1.9673506495862643e-13 K=2.62 tau=9.68044028536725e-08 off=-0.2

*Grain_1004:
XU_1004 in out fe_tanh Vc=0.22754716808666395 Qo=8.023110017000289e-14 K=2.62 tau=8.656959424639174e-08 off=-0.2

*Grain_1005:
XU_1005 in out fe_tanh Vc=0.018485303174196555 Qo=6.517752882237506e-15 K=2.62 tau=1.1309734475319248e-07 off=-0.2

*Grain_1006:
XU_1006 in out fe_tanh Vc=0.6508077510932229 Qo=2.29469003321052e-13 K=2.62 tau=9.300501632136596e-08 off=-0.2

*Grain_1007:
XU_1007 in out fe_tanh Vc=0.7014146913992758 Qo=2.4731255870841637e-13 K=2.62 tau=1.0192637074609956e-07 off=-0.2

*Grain_1008:
XU_1008 in out fe_tanh Vc=0.6312721343268181 Qo=2.225809192422765e-13 K=2.62 tau=1.0833581536886619e-07 off=-0.2

*Grain_1009:
XU_1009 in out fe_tanh Vc=0.7013256066698126 Qo=2.472811482280607e-13 K=2.62 tau=8.847261719812911e-08 off=-0.2

*Grain_1010:
XU_1010 in out fe_tanh Vc=-0.0699612729498646 Qo=2.4667720302823978e-14 K=2.62 tau=1.0134469122657151e-07 off=-0.2

*Grain_1011:
XU_1011 in out fe_tanh Vc=0.7615574667074615 Qo=2.6851836439181317e-13 K=2.62 tau=1.1530514631828598e-07 off=-0.2

*Grain_1012:
XU_1012 in out fe_tanh Vc=0.5297280872899959 Qo=1.86777394733565e-13 K=2.62 tau=9.081218593833672e-08 off=-0.2

*Grain_1013:
XU_1013 in out fe_tanh Vc=0.5827447272794531 Qo=2.0547058871808034e-13 K=2.62 tau=1.1357346968988401e-07 off=-0.2

*Grain_1014:
XU_1014 in out fe_tanh Vc=0.014499081164388916 Qo=5.1122465862991624e-15 K=2.62 tau=9.181020097451606e-08 off=-0.2

*Grain_1015:
XU_1015 in out fe_tanh Vc=0.34025859755463383 Qo=1.1997214403350986e-13 K=2.62 tau=9.750297414236248e-08 off=-0.2

*Grain_1016:
XU_1016 in out fe_tanh Vc=0.22812979662080637 Qo=8.04365297900581e-14 K=2.62 tau=9.055400482604902e-08 off=-0.2

*Grain_1017:
XU_1017 in out fe_tanh Vc=0.5784354392857586 Qo=2.0395117224021046e-13 K=2.62 tau=8.890849485363259e-08 off=-0.2

*Grain_1018:
XU_1018 in out fe_tanh Vc=0.4043229618121948 Qo=1.4256066697271128e-13 K=2.62 tau=1.0618708747045338e-07 off=-0.2

*Grain_1019:
XU_1019 in out fe_tanh Vc=0.5131820610147834 Qo=1.8094341357412256e-13 K=2.62 tau=1.0527058650775883e-07 off=-0.2

*Grain_1020:
XU_1020 in out fe_tanh Vc=0.439684162965204 Qo=1.5502871083233942e-13 K=2.62 tau=1.0542830373474414e-07 off=-0.2

*Grain_1021:
XU_1021 in out fe_tanh Vc=-0.06281731496232729 Qo=2.214882449002221e-14 K=2.62 tau=9.10571421752775e-08 off=-0.2

*Grain_1022:
XU_1022 in out fe_tanh Vc=0.9701628740059627 Qo=3.420707687996586e-13 K=2.62 tau=1.0460742786657289e-07 off=-0.2

*Grain_1023:
XU_1023 in out fe_tanh Vc=-0.14194470546965282 Qo=5.004843601832864e-14 K=2.62 tau=9.37666138932434e-08 off=-0.2

*Grain_1024:
XU_1024 in out fe_tanh Vc=0.345788083129691 Qo=1.2192179128595134e-13 K=2.62 tau=1.198743961682286e-07 off=-0.2

*Grain_1025:
XU_1025 in out fe_tanh Vc=0.9731931141892083 Qo=3.4313920443753286e-13 K=2.62 tau=1.1924230928924768e-07 off=-0.2

*Grain_1026:
XU_1026 in out fe_tanh Vc=0.020455147174567312 Qo=7.212302292111213e-15 K=2.62 tau=1.1915756244765419e-07 off=-0.2

*Grain_1027:
XU_1027 in out fe_tanh Vc=0.5518619309390903 Qo=1.9458159041699066e-13 K=2.62 tau=1.0292059114721778e-07 off=-0.2

*Grain_1028:
XU_1028 in out fe_tanh Vc=0.42022149386061647 Qo=1.4816634744792208e-13 K=2.62 tau=9.519953841396489e-08 off=-0.2

*Grain_1029:
XU_1029 in out fe_tanh Vc=0.8252346584796354 Qo=2.909703737689283e-13 K=2.62 tau=1.0741486385895653e-07 off=-0.2

*Grain_1030:
XU_1030 in out fe_tanh Vc=0.46650251257204156 Qo=1.6448462149821445e-13 K=2.62 tau=1.0851352477751467e-07 off=-0.2

*Grain_1031:
XU_1031 in out fe_tanh Vc=0.09326476406907724 Qo=3.2884323242853706e-14 K=2.62 tau=1.071952035457072e-07 off=-0.2

*Grain_1032:
XU_1032 in out fe_tanh Vc=0.30181455795022094 Qo=1.0641711885619597e-13 K=2.62 tau=1.0449866741633267e-07 off=-0.2

*Grain_1033:
XU_1033 in out fe_tanh Vc=-0.01603207359214187 Qo=5.65276603141069e-15 K=2.62 tau=1.052138654181175e-07 off=-0.2

*Grain_1034:
XU_1034 in out fe_tanh Vc=0.4253186645412935 Qo=1.4996356432784934e-13 K=2.62 tau=1.1506028686206559e-07 off=-0.2

*Grain_1035:
XU_1035 in out fe_tanh Vc=0.5566693423376167 Qo=1.9627664076069205e-13 K=2.62 tau=9.209119879725214e-08 off=-0.2

*Grain_1036:
XU_1036 in out fe_tanh Vc=1.3054755097370265 Qo=4.602990108464265e-13 K=2.62 tau=1.0058810100436996e-07 off=-0.2

*Grain_1037:
XU_1037 in out fe_tanh Vc=0.12957572695860609 Qo=4.5687244612323335e-14 K=2.62 tau=1.009508185248805e-07 off=-0.2

*Grain_1038:
XU_1038 in out fe_tanh Vc=0.7306618389746182 Qo=2.5762484185627983e-13 K=2.62 tau=1.1838224394931767e-07 off=-0.2

*Grain_1039:
XU_1039 in out fe_tanh Vc=0.09556584178032568 Qo=3.369566270228315e-14 K=2.62 tau=8.814715417981332e-08 off=-0.2

*Grain_1040:
XU_1040 in out fe_tanh Vc=0.582076374577052 Qo=2.0523493352155062e-13 K=2.62 tau=1.0714820087487326e-07 off=-0.2

*Grain_1041:
XU_1041 in out fe_tanh Vc=0.019806198864430358 Qo=6.983488911072243e-15 K=2.62 tau=1.0252016342035391e-07 off=-0.2

*Grain_1042:
XU_1042 in out fe_tanh Vc=0.31294220453420685 Qo=1.1034062770600129e-13 K=2.62 tau=1.2331737236891733e-07 off=-0.2

*Grain_1043:
XU_1043 in out fe_tanh Vc=0.6294275481506485 Qo=2.2193053462304846e-13 K=2.62 tau=9.053871983027351e-08 off=-0.2

*Grain_1044:
XU_1044 in out fe_tanh Vc=0.7340838682046127 Qo=2.588314188145648e-13 K=2.62 tau=9.944360811225768e-08 off=-0.2

*Grain_1045:
XU_1045 in out fe_tanh Vc=0.7281443357634976 Qo=2.567371926976104e-13 K=2.62 tau=8.897057241898963e-08 off=-0.2

*Grain_1046:
XU_1046 in out fe_tanh Vc=-0.056460537319967974 Qo=1.9907481439827353e-14 K=2.62 tau=1.199912097847144e-07 off=-0.2

*Grain_1047:
XU_1047 in out fe_tanh Vc=0.7425776047992403 Qo=2.6182623451484916e-13 K=2.62 tau=1.1840321882233686e-07 off=-0.2

*Grain_1048:
XU_1048 in out fe_tanh Vc=0.6619944501365412 Qo=2.3341333354086087e-13 K=2.62 tau=1.0035298135344934e-07 off=-0.2

*Grain_1049:
XU_1049 in out fe_tanh Vc=0.11817886640415715 Qo=4.166881331978668e-14 K=2.62 tau=1.116694574669527e-07 off=-0.2

*Grain_1050:
XU_1050 in out fe_tanh Vc=1.084546598029662 Qo=3.824014487950615e-13 K=2.62 tau=9.788977284246909e-08 off=-0.2

*Grain_1051:
XU_1051 in out fe_tanh Vc=0.8463050672065137 Qo=2.9839961179198827e-13 K=2.62 tau=9.05127324439605e-08 off=-0.2

*Grain_1052:
XU_1052 in out fe_tanh Vc=0.6231128175019915 Qo=2.1970401696748254e-13 K=2.62 tau=1.0662476497158658e-07 off=-0.2

*Grain_1053:
XU_1053 in out fe_tanh Vc=0.6077362753304043 Qo=2.1428238546307712e-13 K=2.62 tau=1.0655588358138639e-07 off=-0.2

*Grain_1054:
XU_1054 in out fe_tanh Vc=1.2029226979236125 Qo=4.2413980488266e-13 K=2.62 tau=1.1516080607215351e-07 off=-0.2

*Grain_1055:
XU_1055 in out fe_tanh Vc=0.02577285980781935 Qo=9.087280295754137e-15 K=2.62 tau=9.520668074347028e-08 off=-0.2

*Grain_1056:
XU_1056 in out fe_tanh Vc=0.2772158853586239 Qo=9.77438464909962e-14 K=2.62 tau=9.840324375988048e-08 off=-0.2

*Grain_1057:
XU_1057 in out fe_tanh Vc=0.025407768811799958 Qo=8.958552469699005e-15 K=2.62 tau=1.1540527686936025e-07 off=-0.2

*Grain_1058:
XU_1058 in out fe_tanh Vc=0.6956691017557597 Qo=2.4528671509058193e-13 K=2.62 tau=9.548083169392996e-08 off=-0.2

*Grain_1059:
XU_1059 in out fe_tanh Vc=0.6320317555822141 Qo=2.2284875491584433e-13 K=2.62 tau=9.199877850750321e-08 off=-0.2

*Grain_1060:
XU_1060 in out fe_tanh Vc=0.01964166911469023 Qo=6.9254771900592265e-15 K=2.62 tau=9.771072708209402e-08 off=-0.2

*Grain_1061:
XU_1061 in out fe_tanh Vc=0.5817530236463911 Qo=2.0512092286993035e-13 K=2.62 tau=1.1185791112866509e-07 off=-0.2

*Grain_1062:
XU_1062 in out fe_tanh Vc=0.8184232955883621 Qo=2.885687480180165e-13 K=2.62 tau=1.0333981601712125e-07 off=-0.2

*Grain_1063:
XU_1063 in out fe_tanh Vc=-0.03909451790190749 Qo=1.3784378018237091e-14 K=2.62 tau=9.976007484712957e-08 off=-0.2

*Grain_1064:
XU_1064 in out fe_tanh Vc=0.7021070821870778 Qo=2.4755668951927214e-13 K=2.62 tau=8.995706544605977e-08 off=-0.2

*Grain_1065:
XU_1065 in out fe_tanh Vc=0.23850042139577726 Qo=8.409311950788448e-14 K=2.62 tau=1.0537012139908986e-07 off=-0.2

*Grain_1066:
XU_1066 in out fe_tanh Vc=0.1265582187020765 Qo=4.4623298138152184e-14 K=2.62 tau=8.782768650047501e-08 off=-0.2

*Grain_1067:
XU_1067 in out fe_tanh Vc=0.6624115077765518 Qo=2.3356038434168476e-13 K=2.62 tau=9.949891491641352e-08 off=-0.2

*Grain_1068:
XU_1068 in out fe_tanh Vc=0.23830708989863938 Qo=8.402495254785015e-14 K=2.62 tau=1.1049657697687592e-07 off=-0.2

*Grain_1069:
XU_1069 in out fe_tanh Vc=0.15723851092668328 Qo=5.544089529576608e-14 K=2.62 tau=1.0400464769600749e-07 off=-0.2

*Grain_1070:
XU_1070 in out fe_tanh Vc=0.6594556121862396 Qo=2.3251816194361e-13 K=2.62 tau=9.765947083910444e-08 off=-0.2

*Grain_1071:
XU_1071 in out fe_tanh Vc=0.32108909575234135 Qo=1.1321314882279815e-13 K=2.62 tau=9.06320716394298e-08 off=-0.2

*Grain_1072:
XU_1072 in out fe_tanh Vc=0.5614725477100289 Qo=1.979702080971325e-13 K=2.62 tau=9.414444031249342e-08 off=-0.2

*Grain_1073:
XU_1073 in out fe_tanh Vc=0.7292657375598462 Qo=2.5713258896032907e-13 K=2.62 tau=9.719049644245585e-08 off=-0.2

*Grain_1074:
XU_1074 in out fe_tanh Vc=0.03403096518490534 Qo=1.1999014532196416e-14 K=2.62 tau=1.0423768899762943e-07 off=-0.2

*Grain_1075:
XU_1075 in out fe_tanh Vc=0.2522450208140383 Qo=8.893934256570373e-14 K=2.62 tau=9.224871750531286e-08 off=-0.2

*Grain_1076:
XU_1076 in out fe_tanh Vc=0.8438815622201403 Qo=2.9754510556824937e-13 K=2.62 tau=9.90720052394489e-08 off=-0.2

*Grain_1077:
XU_1077 in out fe_tanh Vc=0.44097316809685166 Qo=1.5548320253490144e-13 K=2.62 tau=1.2700430161836015e-07 off=-0.2

*Grain_1078:
XU_1078 in out fe_tanh Vc=0.5622740623531891 Qo=1.9825281500524671e-13 K=2.62 tau=8.76523638148339e-08 off=-0.2

*Grain_1079:
XU_1079 in out fe_tanh Vc=-0.18492461076830985 Qo=6.52027669480832e-14 K=2.62 tau=9.790284770372388e-08 off=-0.2

*Grain_1080:
XU_1080 in out fe_tanh Vc=0.8289783384612396 Qo=2.922903619108775e-13 K=2.62 tau=1.026836474086941e-07 off=-0.2

*Grain_1081:
XU_1081 in out fe_tanh Vc=0.6621337578279448 Qo=2.3346245218925996e-13 K=2.62 tau=9.504715771952977e-08 off=-0.2

*Grain_1082:
XU_1082 in out fe_tanh Vc=0.06275715605995869 Qo=2.2127612998081276e-14 K=2.62 tau=1.0440023161791436e-07 off=-0.2

*Grain_1083:
XU_1083 in out fe_tanh Vc=-0.3745169770158618 Qo=1.320513428094266e-13 K=2.62 tau=1.1970871776267226e-07 off=-0.2

*Grain_1084:
XU_1084 in out fe_tanh Vc=0.81780947205686 Qo=2.883523193203678e-13 K=2.62 tau=9.997390708532372e-08 off=-0.2

*Grain_1085:
XU_1085 in out fe_tanh Vc=0.01117312171875634 Qo=3.9395429763720835e-15 K=2.62 tau=9.887758341211871e-08 off=-0.2

*Grain_1086:
XU_1086 in out fe_tanh Vc=0.7145311126764167 Qo=2.5193729176137813e-13 K=2.62 tau=9.572802351931921e-08 off=-0.2

*Grain_1087:
XU_1087 in out fe_tanh Vc=0.478402663029322 Qo=1.6868050831765637e-13 K=2.62 tau=8.76159507305595e-08 off=-0.2

*Grain_1088:
XU_1088 in out fe_tanh Vc=0.02675555028634824 Qo=9.433768186075547e-15 K=2.62 tau=1.1681332779190107e-07 off=-0.2

*Grain_1089:
XU_1089 in out fe_tanh Vc=0.19540127673017937 Qo=6.889674584178791e-14 K=2.62 tau=9.64031320435117e-08 off=-0.2

*Grain_1090:
XU_1090 in out fe_tanh Vc=0.09469686342248235 Qo=3.338926869061547e-14 K=2.62 tau=9.553970652010389e-08 off=-0.2

*Grain_1091:
XU_1091 in out fe_tanh Vc=-0.4610049373839649 Qo=1.6254622556336058e-13 K=2.62 tau=8.306181991269118e-08 off=-0.2

*Grain_1092:
XU_1092 in out fe_tanh Vc=0.7503719894633287 Qo=2.645744649674902e-13 K=2.62 tau=8.433890765944656e-08 off=-0.2

*Grain_1093:
XU_1093 in out fe_tanh Vc=0.3430412175096756 Qo=1.2095327098940756e-13 K=2.62 tau=1.1267311581818099e-07 off=-0.2

*Grain_1094:
XU_1094 in out fe_tanh Vc=0.6557433640756836 Qo=2.312092563988023e-13 K=2.62 tau=1.0329900919507501e-07 off=-0.2

*Grain_1095:
XU_1095 in out fe_tanh Vc=0.4211443485852899 Qo=1.4849173778558355e-13 K=2.62 tau=1.1055267069506763e-07 off=-0.2

*Grain_1096:
XU_1096 in out fe_tanh Vc=1.1248879571491086 Qo=3.9662545189614015e-13 K=2.62 tau=1.0202600351454246e-07 off=-0.2

*Grain_1097:
XU_1097 in out fe_tanh Vc=0.5666082717263448 Qo=1.9978101853904316e-13 K=2.62 tau=9.422806280731106e-08 off=-0.2

*Grain_1098:
XU_1098 in out fe_tanh Vc=0.17001899424135353 Qo=5.994717962205498e-14 K=2.62 tau=9.293958094527789e-08 off=-0.2

*Grain_1099:
XU_1099 in out fe_tanh Vc=0.3075107057615492 Qo=1.084255297253647e-13 K=2.62 tau=1.0029007835685794e-07 off=-0.2

*Grain_1100:
XU_1100 in out fe_tanh Vc=-0.03913108664798104 Qo=1.3797271831656034e-14 K=2.62 tau=1.087089157447349e-07 off=-0.2

*Grain_1101:
XU_1101 in out fe_tanh Vc=0.5998066183601215 Qo=2.114864592028381e-13 K=2.62 tau=1.0265244330145215e-07 off=-0.2

*Grain_1102:
XU_1102 in out fe_tanh Vc=0.49216085080830124 Qo=1.7353152251016254e-13 K=2.62 tau=1.1666554292924047e-07 off=-0.2

*Grain_1103:
XU_1103 in out fe_tanh Vc=0.6575156201296233 Qo=2.318341380626179e-13 K=2.62 tau=1.0647773297980678e-07 off=-0.2

*Grain_1104:
XU_1104 in out fe_tanh Vc=0.6974164894412294 Qo=2.4590282838967317e-13 K=2.62 tau=1.1113360043098541e-07 off=-0.2

*Grain_1105:
XU_1105 in out fe_tanh Vc=0.4114200099717905 Qo=1.4506302279894155e-13 K=2.62 tau=1.1380405189445324e-07 off=-0.2

*Grain_1106:
XU_1106 in out fe_tanh Vc=0.2318541797732146 Qo=8.174971404229423e-14 K=2.62 tau=1.0596638405261644e-07 off=-0.2

*Grain_1107:
XU_1107 in out fe_tanh Vc=0.41734415137627134 Qo=1.471518221737733e-13 K=2.62 tau=9.478187497689827e-08 off=-0.2

*Grain_1108:
XU_1108 in out fe_tanh Vc=0.45793510478376337 Qo=1.6146382999270639e-13 K=2.62 tau=9.41731237169699e-08 off=-0.2

*Grain_1109:
XU_1109 in out fe_tanh Vc=0.47416853286382293 Qo=1.6718759181907968e-13 K=2.62 tau=9.660605581511685e-08 off=-0.2

*Grain_1110:
XU_1110 in out fe_tanh Vc=0.8527167845343016 Qo=3.006603260848226e-13 K=2.62 tau=1.0166687468166762e-07 off=-0.2

*Grain_1111:
XU_1111 in out fe_tanh Vc=0.42860374499159665 Qo=1.5112185436894716e-13 K=2.62 tau=1.0402519831070774e-07 off=-0.2

*Grain_1112:
XU_1112 in out fe_tanh Vc=0.3156606496698954 Qo=1.1129912719347904e-13 K=2.62 tau=9.164516695760817e-08 off=-0.2

*Grain_1113:
XU_1113 in out fe_tanh Vc=0.31102951737015494 Qo=1.096662312863786e-13 K=2.62 tau=9.633154446343784e-08 off=-0.2

*Grain_1114:
XU_1114 in out fe_tanh Vc=0.7985990733381488 Qo=2.8157890422201064e-13 K=2.62 tau=1.0110180646166746e-07 off=-0.2

*Grain_1115:
XU_1115 in out fe_tanh Vc=0.700497470637716 Qo=2.4698915485585474e-13 K=2.62 tau=8.219953295734467e-08 off=-0.2

*Grain_1116:
XU_1116 in out fe_tanh Vc=0.5328317186778638 Qo=1.8787170745503101e-13 K=2.62 tau=1.0171290570211645e-07 off=-0.2

*Grain_1117:
XU_1117 in out fe_tanh Vc=0.3913498829745643 Qo=1.379864751843131e-13 K=2.62 tau=1.0962351464485046e-07 off=-0.2

*Grain_1118:
XU_1118 in out fe_tanh Vc=0.13065601040412028 Qo=4.6068142911598296e-14 K=2.62 tau=1.1547122205826525e-07 off=-0.2

*Grain_1119:
XU_1119 in out fe_tanh Vc=0.5600149611668599 Qo=1.9745627609378237e-13 K=2.62 tau=8.888343813174927e-08 off=-0.2

*Grain_1120:
XU_1120 in out fe_tanh Vc=0.6321724406762406 Qo=2.2289835922411224e-13 K=2.62 tau=1.0130382749741734e-07 off=-0.2

*Grain_1121:
XU_1121 in out fe_tanh Vc=0.665022387402586 Qo=2.3448095719068805e-13 K=2.62 tau=8.677001379750975e-08 off=-0.2

*Grain_1122:
XU_1122 in out fe_tanh Vc=0.34438383227743957 Qo=1.2142666497109478e-13 K=2.62 tau=1.1640917841742619e-07 off=-0.2

*Grain_1123:
XU_1123 in out fe_tanh Vc=0.4881379731430048 Qo=1.7211309175732128e-13 K=2.62 tau=1.0722870523188304e-07 off=-0.2

*Grain_1124:
XU_1124 in out fe_tanh Vc=0.32003798567792424 Qo=1.1284253679374341e-13 K=2.62 tau=9.066458615907727e-08 off=-0.2

*Grain_1125:
XU_1125 in out fe_tanh Vc=0.4330730546372831 Qo=1.5269769305280746e-13 K=2.62 tau=1.0126707870657564e-07 off=-0.2

*Grain_1126:
XU_1126 in out fe_tanh Vc=0.39956351998111733 Qo=1.4088253027027143e-13 K=2.62 tau=1.0692725025176374e-07 off=-0.2

*Grain_1127:
XU_1127 in out fe_tanh Vc=0.3697285444301011 Qo=1.3036298422568387e-13 K=2.62 tau=1.0703700789970743e-07 off=-0.2

*Grain_1128:
XU_1128 in out fe_tanh Vc=0.9790348918288976 Qo=3.451989630841546e-13 K=2.62 tau=9.253660187167164e-08 off=-0.2

*Grain_1129:
XU_1129 in out fe_tanh Vc=0.4147839972764127 Qo=1.4624913469247636e-13 K=2.62 tau=1.0556373355510372e-07 off=-0.2

*Grain_1130:
XU_1130 in out fe_tanh Vc=0.34879541933987585 Qo=1.2298215118738644e-13 K=2.62 tau=9.54524072670435e-08 off=-0.2

*Grain_1131:
XU_1131 in out fe_tanh Vc=0.9240669433914048 Qo=3.258177551600534e-13 K=2.62 tau=7.342480309258378e-08 off=-0.2

*Grain_1132:
XU_1132 in out fe_tanh Vc=0.37344290326194984 Qo=1.3167263399197712e-13 K=2.62 tau=9.92411019378071e-08 off=-0.2

*Grain_1133:
XU_1133 in out fe_tanh Vc=1.0878280566880711 Qo=3.83558461824669e-13 K=2.62 tau=9.456197132769797e-08 off=-0.2

*Grain_1134:
XU_1134 in out fe_tanh Vc=0.2764505769127211 Qo=9.747400556482485e-14 K=2.62 tau=1.0964546566200876e-07 off=-0.2

*Grain_1135:
XU_1135 in out fe_tanh Vc=0.7917897308130953 Qo=2.7917799083419226e-13 K=2.62 tau=9.6334435891904e-08 off=-0.2

*Grain_1136:
XU_1136 in out fe_tanh Vc=0.30036246718188053 Qo=1.0590512461398996e-13 K=2.62 tau=9.866160051196162e-08 off=-0.2

*Grain_1137:
XU_1137 in out fe_tanh Vc=0.6392919006206175 Qo=2.2540861724558794e-13 K=2.62 tau=8.168342357928457e-08 off=-0.2

*Grain_1138:
XU_1138 in out fe_tanh Vc=0.359013876372991 Qo=1.2658508791782507e-13 K=2.62 tau=9.53958051854656e-08 off=-0.2

*Grain_1139:
XU_1139 in out fe_tanh Vc=0.6138001031580598 Qo=2.1642043702374953e-13 K=2.62 tau=9.206017345943617e-08 off=-0.2

*Grain_1140:
XU_1140 in out fe_tanh Vc=0.6163354810814232 Qo=2.1731438864638942e-13 K=2.62 tau=1.082491997568067e-07 off=-0.2

*Grain_1141:
XU_1141 in out fe_tanh Vc=0.5660923184631442 Qo=1.9959909802431668e-13 K=2.62 tau=9.678970256885584e-08 off=-0.2

*Grain_1142:
XU_1142 in out fe_tanh Vc=0.4527611136777363 Qo=1.5963952691657116e-13 K=2.62 tau=1.0443310452362257e-07 off=-0.2

*Grain_1143:
XU_1143 in out fe_tanh Vc=0.5390806137591605 Qo=1.900750120772551e-13 K=2.62 tau=8.814119050375038e-08 off=-0.2

*Grain_1144:
XU_1144 in out fe_tanh Vc=0.28522609948449684 Qo=1.0056817648516831e-13 K=2.62 tau=9.179036855218889e-08 off=-0.2

*Grain_1145:
XU_1145 in out fe_tanh Vc=0.47868160183563024 Qo=1.6877885965069382e-13 K=2.62 tau=1.0371457580837307e-07 off=-0.2

*Grain_1146:
XU_1146 in out fe_tanh Vc=0.37263543308322356 Qo=1.3138792721518698e-13 K=2.62 tau=1.0402417499091644e-07 off=-0.2

*Grain_1147:
XU_1147 in out fe_tanh Vc=0.12099185960626324 Qo=4.2660649611459424e-14 K=2.62 tau=9.47281566991971e-08 off=-0.2

*Grain_1148:
XU_1148 in out fe_tanh Vc=0.13891676119158558 Qo=4.898080989612493e-14 K=2.62 tau=8.87151280702035e-08 off=-0.2

*Grain_1149:
XU_1149 in out fe_tanh Vc=0.07631987621640735 Qo=2.6909707051808694e-14 K=2.62 tau=1.202464154351341e-07 off=-0.2

*Grain_1150:
XU_1150 in out fe_tanh Vc=0.5945603745454888 Qo=2.0963668046664333e-13 K=2.62 tau=9.378100999049545e-08 off=-0.2

*Grain_1151:
XU_1151 in out fe_tanh Vc=0.41496863143671747 Qo=1.4631423504918383e-13 K=2.62 tau=9.087696573648405e-08 off=-0.2

*Grain_1152:
XU_1152 in out fe_tanh Vc=0.35082389561218397 Qo=1.2369737381293917e-13 K=2.62 tau=1.022010561906786e-07 off=-0.2

*Grain_1153:
XU_1153 in out fe_tanh Vc=0.5860199468686591 Qo=2.0662540190758246e-13 K=2.62 tau=9.614103705919891e-08 off=-0.2

*Grain_1154:
XU_1154 in out fe_tanh Vc=0.6633212808790347 Qo=2.338811622161406e-13 K=2.62 tau=9.355744049260318e-08 off=-0.2

*Grain_1155:
XU_1155 in out fe_tanh Vc=0.5897161199902505 Qo=2.0792863955478154e-13 K=2.62 tau=1.1000161373923099e-07 off=-0.2

*Grain_1156:
XU_1156 in out fe_tanh Vc=0.9243343326258582 Qo=3.25912034217157e-13 K=2.62 tau=1.15642477055192e-07 off=-0.2

*Grain_1157:
XU_1157 in out fe_tanh Vc=1.269308376534352 Qo=4.4754680254058434e-13 K=2.62 tau=1.0323358986648493e-07 off=-0.2

*Grain_1158:
XU_1158 in out fe_tanh Vc=0.3240617562568405 Qo=1.1426128237995605e-13 K=2.62 tau=9.646857304407577e-08 off=-0.2

*Grain_1159:
XU_1159 in out fe_tanh Vc=0.27599813320795274 Qo=9.731447795345623e-14 K=2.62 tau=1.0790477367233102e-07 off=-0.2

*Grain_1160:
XU_1160 in out fe_tanh Vc=0.08924270433381387 Qo=3.14661808848405e-14 K=2.62 tau=1.1155938681419938e-07 off=-0.2

*Grain_1161:
XU_1161 in out fe_tanh Vc=0.9312638560015015 Qo=3.283553223000475e-13 K=2.62 tau=1.0461210736997101e-07 off=-0.2

*Grain_1162:
XU_1162 in out fe_tanh Vc=0.6743517715241664 Qo=2.3777041474921e-13 K=2.62 tau=9.297606685404294e-08 off=-0.2

*Grain_1163:
XU_1163 in out fe_tanh Vc=0.7405508222260193 Qo=2.61111609072475e-13 K=2.62 tau=8.991964449644739e-08 off=-0.2

*Grain_1164:
XU_1164 in out fe_tanh Vc=0.22722215084515585 Qo=8.011650199205289e-14 K=2.62 tau=9.139503410947914e-08 off=-0.2

*Grain_1165:
XU_1165 in out fe_tanh Vc=0.3387326261769785 Qo=1.1943410014798636e-13 K=2.62 tau=1.1617522047573822e-07 off=-0.2

*Grain_1166:
XU_1166 in out fe_tanh Vc=0.3600363722840997 Qo=1.2694561084833385e-13 K=2.62 tau=9.410939375779756e-08 off=-0.2

*Grain_1167:
XU_1167 in out fe_tanh Vc=0.4184446358140172 Qo=1.4753984316257634e-13 K=2.62 tau=1.015867076928529e-07 off=-0.2

*Grain_1168:
XU_1168 in out fe_tanh Vc=0.343799357680886 Qo=1.2122058444591304e-13 K=2.62 tau=1.1417452842578043e-07 off=-0.2

*Grain_1169:
XU_1169 in out fe_tanh Vc=0.6522572998245594 Qo=2.2998010126370307e-13 K=2.62 tau=1.0636676462382074e-07 off=-0.2

*Grain_1170:
XU_1170 in out fe_tanh Vc=0.5040064397798697 Qo=1.7770817143680893e-13 K=2.62 tau=1.2038457036125056e-07 off=-0.2

*Grain_1171:
XU_1171 in out fe_tanh Vc=0.6804096830272086 Qo=2.399063802666384e-13 K=2.62 tau=9.765116599737465e-08 off=-0.2

*Grain_1172:
XU_1172 in out fe_tanh Vc=0.4951215530255732 Qo=1.7457543968199493e-13 K=2.62 tau=9.800363827198431e-08 off=-0.2

*Grain_1173:
XU_1173 in out fe_tanh Vc=1.0531965895414432 Qo=3.713477156614074e-13 K=2.62 tau=9.460056585922539e-08 off=-0.2

*Grain_1174:
XU_1174 in out fe_tanh Vc=0.9046141034492874 Qo=3.1895885745057883e-13 K=2.62 tau=1.1237441300612687e-07 off=-0.2

*Grain_1175:
XU_1175 in out fe_tanh Vc=0.38198167525874627 Qo=1.346833287730384e-13 K=2.62 tau=8.231394692873353e-08 off=-0.2

*Grain_1176:
XU_1176 in out fe_tanh Vc=0.03880752870166343 Qo=1.3683188188163175e-14 K=2.62 tau=8.385715355242357e-08 off=-0.2

*Grain_1177:
XU_1177 in out fe_tanh Vc=0.11188465593698627 Qo=3.944953089703055e-14 K=2.62 tau=8.096601990059329e-08 off=-0.2

*Grain_1178:
XU_1178 in out fe_tanh Vc=0.5393845448066849 Qo=1.901821754514414e-13 K=2.62 tau=9.422588893027024e-08 off=-0.2

*Grain_1179:
XU_1179 in out fe_tanh Vc=1.1755156958107336 Qo=4.1447634059801376e-13 K=2.62 tau=9.873414967920903e-08 off=-0.2

*Grain_1180:
XU_1180 in out fe_tanh Vc=1.0641963548735414 Qo=3.752261347233839e-13 K=2.62 tau=1.1004710975247214e-07 off=-0.2

*Grain_1181:
XU_1181 in out fe_tanh Vc=0.7148484716081978 Qo=2.520491896876836e-13 K=2.62 tau=1.163700229675871e-07 off=-0.2

*Grain_1182:
XU_1182 in out fe_tanh Vc=0.5987369926386246 Qo=2.111093187219109e-13 K=2.62 tau=1.2259118445393093e-07 off=-0.2

*Grain_1183:
XU_1183 in out fe_tanh Vc=0.7815059684127619 Qo=2.7555202801424886e-13 K=2.62 tau=1.0684321494356015e-07 off=-0.2

*Grain_1184:
XU_1184 in out fe_tanh Vc=0.642300658186425 Qo=2.2646947830432726e-13 K=2.62 tau=1.0341986145507964e-07 off=-0.2

*Grain_1185:
XU_1185 in out fe_tanh Vc=0.16558189137227147 Qo=5.838269676011777e-14 K=2.62 tau=1.0761748760927593e-07 off=-0.2

*Grain_1186:
XU_1186 in out fe_tanh Vc=0.8595131006281864 Qo=3.0305664646929695e-13 K=2.62 tau=9.442670040372047e-08 off=-0.2

*Grain_1187:
XU_1187 in out fe_tanh Vc=0.5031188828934055 Qo=1.7739522680179872e-13 K=2.62 tau=1.016375292120734e-07 off=-0.2

*Grain_1188:
XU_1188 in out fe_tanh Vc=0.5595819598566588 Qo=1.9730360369717729e-13 K=2.62 tau=1.0941586605120168e-07 off=-0.2

*Grain_1189:
XU_1189 in out fe_tanh Vc=0.748470057719669 Qo=2.6390386081308497e-13 K=2.62 tau=1.1405744618990004e-07 off=-0.2

*Grain_1190:
XU_1190 in out fe_tanh Vc=0.8981383814674933 Qo=3.1667557568810687e-13 K=2.62 tau=9.319204053604061e-08 off=-0.2

*Grain_1191:
XU_1191 in out fe_tanh Vc=0.07524020061075831 Qo=2.652902307144404e-14 K=2.62 tau=9.06245066200697e-08 off=-0.2

*Grain_1192:
XU_1192 in out fe_tanh Vc=0.3773365040261838 Qo=1.3304548286354946e-13 K=2.62 tau=9.585031581842783e-08 off=-0.2

*Grain_1193:
XU_1193 in out fe_tanh Vc=0.907959658498636 Qo=3.201384702954476e-13 K=2.62 tau=8.863161418893279e-08 off=-0.2

*Grain_1194:
XU_1194 in out fe_tanh Vc=0.49827184706130534 Qo=1.7568620523654372e-13 K=2.62 tau=1.1139791602309342e-07 off=-0.2

*Grain_1195:
XU_1195 in out fe_tanh Vc=0.8000975418735612 Qo=2.8210725085087524e-13 K=2.62 tau=1.0471898594061603e-07 off=-0.2

*Grain_1196:
XU_1196 in out fe_tanh Vc=-0.09807865758733975 Qo=3.458165912410866e-14 K=2.62 tau=1.0478748613993894e-07 off=-0.2

*Grain_1197:
XU_1197 in out fe_tanh Vc=0.7211696229090809 Qo=2.5427797120790776e-13 K=2.62 tau=1.0590336137773363e-07 off=-0.2

*Grain_1198:
XU_1198 in out fe_tanh Vc=-0.1325656855681538 Qo=4.6741477326902404e-14 K=2.62 tau=9.499735526363866e-08 off=-0.2

*Grain_1199:
XU_1199 in out fe_tanh Vc=0.6368584623120862 Qo=2.2455060862113017e-13 K=2.62 tau=9.776968927558772e-08 off=-0.2

*Grain_1200:
XU_1200 in out fe_tanh Vc=0.5273336238372918 Qo=1.8593312829534613e-13 K=2.62 tau=9.405415426391757e-08 off=-0.2

*Grain_1201:
XU_1201 in out fe_tanh Vc=0.3275248475083216 Qo=1.1548233744045944e-13 K=2.62 tau=8.554201903224125e-08 off=-0.2

*Grain_1202:
XU_1202 in out fe_tanh Vc=0.22566732617584478 Qo=7.956828469346283e-14 K=2.62 tau=8.069945001213043e-08 off=-0.2

*Grain_1203:
XU_1203 in out fe_tanh Vc=0.8146952806994932 Qo=2.872542832479245e-13 K=2.62 tau=1.1277430508449616e-07 off=-0.2

*Grain_1204:
XU_1204 in out fe_tanh Vc=0.8230428534741854 Qo=2.901975628900937e-13 K=2.62 tau=8.477430191614321e-08 off=-0.2

*Grain_1205:
XU_1205 in out fe_tanh Vc=0.3098205650582138 Qo=1.0923996549341929e-13 K=2.62 tau=9.553876946947932e-08 off=-0.2

*Grain_1206:
XU_1206 in out fe_tanh Vc=0.45075431725218446 Qo=1.5893194841145025e-13 K=2.62 tau=1.0933352799252439e-07 off=-0.2

*Grain_1207:
XU_1207 in out fe_tanh Vc=0.5416318062178851 Qo=1.909745397638881e-13 K=2.62 tau=1.0435656818321661e-07 off=-0.2

*Grain_1208:
XU_1208 in out fe_tanh Vc=-0.004843510223610903 Qo=1.7077784671745799e-15 K=2.62 tau=1.1617981424599559e-07 off=-0.2

*Grain_1209:
XU_1209 in out fe_tanh Vc=0.4604693366898786 Qo=1.6235737753989495e-13 K=2.62 tau=9.219015782937414e-08 off=-0.2

*Grain_1210:
XU_1210 in out fe_tanh Vc=0.957482549151708 Qo=3.3759979945240485e-13 K=2.62 tau=1.0232538286160706e-07 off=-0.2

*Grain_1211:
XU_1211 in out fe_tanh Vc=0.6073347240944393 Qo=2.1414080208189518e-13 K=2.62 tau=9.175594297402151e-08 off=-0.2

*Grain_1212:
XU_1212 in out fe_tanh Vc=0.13262517523098805 Qo=4.6762452850957784e-14 K=2.62 tau=9.508424600466333e-08 off=-0.2

*Grain_1213:
XU_1213 in out fe_tanh Vc=0.7467201470007125 Qo=2.6328685791490923e-13 K=2.62 tau=9.60897529586376e-08 off=-0.2

*Grain_1214:
XU_1214 in out fe_tanh Vc=0.6811653049676194 Qo=2.4017280581744404e-13 K=2.62 tau=8.052354040133906e-08 off=-0.2

*Grain_1215:
XU_1215 in out fe_tanh Vc=0.4882633023302122 Qo=1.721572817099259e-13 K=2.62 tau=9.841937906694545e-08 off=-0.2

*Grain_1216:
XU_1216 in out fe_tanh Vc=0.2905135615566855 Qo=1.0243248841102489e-13 K=2.62 tau=1.143417997839898e-07 off=-0.2

*Grain_1217:
XU_1217 in out fe_tanh Vc=0.6958924880639797 Qo=2.4536547910870663e-13 K=2.62 tau=1.167962966773556e-07 off=-0.2

*Grain_1218:
XU_1218 in out fe_tanh Vc=0.6408190863359431 Qo=2.259470892957337e-13 K=2.62 tau=1.1544471779638569e-07 off=-0.2

*Grain_1219:
XU_1219 in out fe_tanh Vc=0.3263161381888875 Qo=1.1505615732448895e-13 K=2.62 tau=9.714162000664767e-08 off=-0.2

*Grain_1220:
XU_1220 in out fe_tanh Vc=0.6525412477636217 Qo=2.300802187722334e-13 K=2.62 tau=1.0024217726070664e-07 off=-0.2

*Grain_1221:
XU_1221 in out fe_tanh Vc=0.5237252385122199 Qo=1.8466084384152445e-13 K=2.62 tau=9.646576902105979e-08 off=-0.2

*Grain_1222:
XU_1222 in out fe_tanh Vc=0.4629058844498176 Qo=1.6321648252916123e-13 K=2.62 tau=1.0895095391074099e-07 off=-0.2

*Grain_1223:
XU_1223 in out fe_tanh Vc=0.36789033502488205 Qo=1.2971484799896801e-13 K=2.62 tau=9.682372942565692e-08 off=-0.2

*Grain_1224:
XU_1224 in out fe_tanh Vc=0.38294059966845684 Qo=1.3502143695965248e-13 K=2.62 tau=9.739310138380703e-08 off=-0.2

*Grain_1225:
XU_1225 in out fe_tanh Vc=0.9191305067275948 Qo=3.240772116596123e-13 K=2.62 tau=1.0617555662121758e-07 off=-0.2

*Grain_1226:
XU_1226 in out fe_tanh Vc=0.4585502884374101 Qo=1.6168073825728155e-13 K=2.62 tau=1.1061297149758002e-07 off=-0.2

*Grain_1227:
XU_1227 in out fe_tanh Vc=0.6731241149192791 Qo=2.3733755398952983e-13 K=2.62 tau=1.028120382189042e-07 off=-0.2

*Grain_1228:
XU_1228 in out fe_tanh Vc=0.1895201033876105 Qo=6.682309662201346e-14 K=2.62 tau=9.878698267483231e-08 off=-0.2

*Grain_1229:
XU_1229 in out fe_tanh Vc=0.7027775689475033 Qo=2.477930971656106e-13 K=2.62 tau=1.1219501343482493e-07 off=-0.2

*Grain_1230:
XU_1230 in out fe_tanh Vc=0.2719113972801004 Qo=9.58735313472959e-14 K=2.62 tau=1.0119530525988029e-07 off=-0.2

*Grain_1231:
XU_1231 in out fe_tanh Vc=0.5407480540135281 Qo=1.906629366258248e-13 K=2.62 tau=1.0655306063258541e-07 off=-0.2

*Grain_1232:
XU_1232 in out fe_tanh Vc=0.4316230381077077 Qo=1.521864301686734e-13 K=2.62 tau=8.693719836018439e-08 off=-0.2

*Grain_1233:
XU_1233 in out fe_tanh Vc=0.7226295521217871 Qo=2.5479272921562393e-13 K=2.62 tau=1.1015268838535675e-07 off=-0.2

*Grain_1234:
XU_1234 in out fe_tanh Vc=-0.058563420746578 Qo=2.0648939363759545e-14 K=2.62 tau=1.1162166628267046e-07 off=-0.2

*Grain_1235:
XU_1235 in out fe_tanh Vc=-0.14894635789840244 Qo=5.251715616145345e-14 K=2.62 tau=1.0358887006529165e-07 off=-0.2

*Grain_1236:
XU_1236 in out fe_tanh Vc=0.5213589181500285 Qo=1.8382650040578905e-13 K=2.62 tau=9.60093296794216e-08 off=-0.2

*Grain_1237:
XU_1237 in out fe_tanh Vc=0.5574804096196903 Qo=1.9656261584401138e-13 K=2.62 tau=1.0933511586797744e-07 off=-0.2

*Grain_1238:
XU_1238 in out fe_tanh Vc=0.27241779822341894 Qo=9.60520837993049e-14 K=2.62 tau=1.0184605855141938e-07 off=-0.2

*Grain_1239:
XU_1239 in out fe_tanh Vc=0.2930958180532369 Qo=1.0334296900008918e-13 K=2.62 tau=1.0577350754234517e-07 off=-0.2

*Grain_1240:
XU_1240 in out fe_tanh Vc=-0.2476844024339359 Qo=8.733130923719493e-14 K=2.62 tau=9.278796287732511e-08 off=-0.2

*Grain_1241:
XU_1241 in out fe_tanh Vc=0.8346338231755831 Qo=2.9428443533504596e-13 K=2.62 tau=1.0837215825603513e-07 off=-0.2

*Grain_1242:
XU_1242 in out fe_tanh Vc=0.780448134010052 Qo=2.751790450470657e-13 K=2.62 tau=9.343945360703371e-08 off=-0.2

*Grain_1243:
XU_1243 in out fe_tanh Vc=0.43398014158622633 Qo=1.530175238135043e-13 K=2.62 tau=1.026353195543541e-07 off=-0.2

*Grain_1244:
XU_1244 in out fe_tanh Vc=-0.023463291867157787 Qo=8.272947257225299e-15 K=2.62 tau=1.1181270353253684e-07 off=-0.2

*Grain_1245:
XU_1245 in out fe_tanh Vc=0.5160582505796492 Qo=1.8195753233915496e-13 K=2.62 tau=1.0684188404524959e-07 off=-0.2

*Grain_1246:
XU_1246 in out fe_tanh Vc=0.32093943239481404 Qo=1.1316037885896815e-13 K=2.62 tau=9.779637197363501e-08 off=-0.2

*Grain_1247:
XU_1247 in out fe_tanh Vc=0.8539293004448365 Qo=3.0108784837083406e-13 K=2.62 tau=9.150405920883843e-08 off=-0.2

*Grain_1248:
XU_1248 in out fe_tanh Vc=0.15287297679906015 Qo=5.390164693317824e-14 K=2.62 tau=1.032430867220279e-07 off=-0.2

*Grain_1249:
XU_1249 in out fe_tanh Vc=0.14757762054086676 Qo=5.203455158780723e-14 K=2.62 tau=9.907213917634755e-08 off=-0.2

*Grain_1250:
XU_1250 in out fe_tanh Vc=0.4135085726430833 Qo=1.4579943135238924e-13 K=2.62 tau=1.0186703412985043e-07 off=-0.2

*Grain_1251:
XU_1251 in out fe_tanh Vc=0.37495148223531266 Qo=1.3220454547100786e-13 K=2.62 tau=9.35662386372694e-08 off=-0.2

*Grain_1252:
XU_1252 in out fe_tanh Vc=0.6307494087244903 Qo=2.2239661086122993e-13 K=2.62 tau=1.1530858406304813e-07 off=-0.2

*Grain_1253:
XU_1253 in out fe_tanh Vc=0.2671740310068261 Qo=9.420317828947053e-14 K=2.62 tau=9.934060764206194e-08 off=-0.2

*Grain_1254:
XU_1254 in out fe_tanh Vc=0.2231098340680932 Qo=7.866653580681944e-14 K=2.62 tau=1.0979030275786355e-07 off=-0.2

*Grain_1255:
XU_1255 in out fe_tanh Vc=0.0780656022397147 Qo=2.7525234463655055e-14 K=2.62 tau=1.0129490904625799e-07 off=-0.2

*Grain_1256:
XU_1256 in out fe_tanh Vc=0.7253634784509342 Qo=2.5575668723371567e-13 K=2.62 tau=9.227849490507391e-08 off=-0.2

*Grain_1257:
XU_1257 in out fe_tanh Vc=0.27144089335026567 Qo=9.570763586179124e-14 K=2.62 tau=9.154820900908028e-08 off=-0.2

*Grain_1258:
XU_1258 in out fe_tanh Vc=0.44093540963021927 Qo=1.55469889236634e-13 K=2.62 tau=9.77906242114762e-08 off=-0.2

*Grain_1259:
XU_1259 in out fe_tanh Vc=0.6383064318700018 Qo=2.2506114976133016e-13 K=2.62 tau=1.0849975700133816e-07 off=-0.2

*Grain_1260:
XU_1260 in out fe_tanh Vc=0.7474039083971762 Qo=2.6352794607941307e-13 K=2.62 tau=9.822625484373415e-08 off=-0.2

*Grain_1261:
XU_1261 in out fe_tanh Vc=0.8062197605471473 Qo=2.8426589050257183e-13 K=2.62 tau=9.839878459850104e-08 off=-0.2

*Grain_1262:
XU_1262 in out fe_tanh Vc=0.43722706293748625 Qo=1.54162359296923e-13 K=2.62 tau=9.000222712016601e-08 off=-0.2

*Grain_1263:
XU_1263 in out fe_tanh Vc=0.12463305921378337 Qo=4.3944504088341595e-14 K=2.62 tau=1.0913417922645032e-07 off=-0.2

*Grain_1264:
XU_1264 in out fe_tanh Vc=0.5652079542714598 Qo=1.9928727910498486e-13 K=2.62 tau=1.1114247646696157e-07 off=-0.2

*Grain_1265:
XU_1265 in out fe_tanh Vc=0.16370293309819473 Qo=5.772019284600494e-14 K=2.62 tau=1.1009095329521173e-07 off=-0.2

*Grain_1266:
XU_1266 in out fe_tanh Vc=0.22058969502678719 Qo=7.777795727795657e-14 K=2.62 tau=9.292697610851863e-08 off=-0.2

*Grain_1267:
XU_1267 in out fe_tanh Vc=0.5671642966052101 Qo=1.9997706794773663e-13 K=2.62 tau=8.629670401446417e-08 off=-0.2

*Grain_1268:
XU_1268 in out fe_tanh Vc=0.6039849145825524 Qo=2.1295968915151464e-13 K=2.62 tau=1.085750345940733e-07 off=-0.2

*Grain_1269:
XU_1269 in out fe_tanh Vc=0.4735833634115933 Qo=1.669812662939895e-13 K=2.62 tau=1.0513324152308027e-07 off=-0.2

*Grain_1270:
XU_1270 in out fe_tanh Vc=0.7656521714462217 Qo=2.6996212072956256e-13 K=2.62 tau=1.006522505325744e-07 off=-0.2

*Grain_1271:
XU_1271 in out fe_tanh Vc=0.3493091432499186 Qo=1.2316328565209079e-13 K=2.62 tau=9.519912863991038e-08 off=-0.2

*Grain_1272:
XU_1272 in out fe_tanh Vc=0.8134255293921828 Qo=2.868065802719464e-13 K=2.62 tau=1.055511591852481e-07 off=-0.2

*Grain_1273:
XU_1273 in out fe_tanh Vc=0.07281415457417628 Qo=2.567362089608531e-14 K=2.62 tau=1.1075156669299761e-07 off=-0.2

*Grain_1274:
XU_1274 in out fe_tanh Vc=0.31889304985628464 Qo=1.1243884264379377e-13 K=2.62 tau=1.2018630585052803e-07 off=-0.2

*Grain_1275:
XU_1275 in out fe_tanh Vc=0.22493623416859512 Qo=7.931050817811287e-14 K=2.62 tau=9.602445740688599e-08 off=-0.2

*Grain_1276:
XU_1276 in out fe_tanh Vc=0.33292092899127657 Qo=1.1738494760091448e-13 K=2.62 tau=1.161026914623464e-07 off=-0.2

*Grain_1277:
XU_1277 in out fe_tanh Vc=0.5369534093980837 Qo=1.8932497880894116e-13 K=2.62 tau=1.1056474925231077e-07 off=-0.2

*Grain_1278:
XU_1278 in out fe_tanh Vc=0.3869161762480016 Qo=1.364231897719111e-13 K=2.62 tau=9.731635698184378e-08 off=-0.2

*Grain_1279:
XU_1279 in out fe_tanh Vc=0.5955101446255533 Qo=2.0997156091834424e-13 K=2.62 tau=1.1846279649254583e-07 off=-0.2

*Grain_1280:
XU_1280 in out fe_tanh Vc=0.5283477355698748 Qo=1.8629069503935173e-13 K=2.62 tau=8.695976670889014e-08 off=-0.2

*Grain_1281:
XU_1281 in out fe_tanh Vc=0.2505448391243461 Qo=8.833987367931906e-14 K=2.62 tau=1.0009938092654871e-07 off=-0.2

*Grain_1282:
XU_1282 in out fe_tanh Vc=0.5465095363589547 Qo=1.9269438386847988e-13 K=2.62 tau=1.1101283068592839e-07 off=-0.2

*Grain_1283:
XU_1283 in out fe_tanh Vc=0.2509500869730751 Qo=8.848276045316222e-14 K=2.62 tau=8.415553688512635e-08 off=-0.2

*Grain_1284:
XU_1284 in out fe_tanh Vc=0.5734282711345045 Qo=2.0218568944871156e-13 K=2.62 tau=9.714438681706455e-08 off=-0.2

*Grain_1285:
XU_1285 in out fe_tanh Vc=0.7484974002443039 Qo=2.6391350154318645e-13 K=2.62 tau=1.0149237674987535e-07 off=-0.2

*Grain_1286:
XU_1286 in out fe_tanh Vc=0.6758063135628454 Qo=2.382832732874551e-13 K=2.62 tau=8.727162651904842e-08 off=-0.2

*Grain_1287:
XU_1287 in out fe_tanh Vc=-0.07005534251320006 Qo=2.4700888391103772e-14 K=2.62 tau=1.0413325909587313e-07 off=-0.2

*Grain_1288:
XU_1288 in out fe_tanh Vc=0.26653587276744206 Qo=9.397816939105684e-14 K=2.62 tau=1.0848133127134597e-07 off=-0.2

*Grain_1289:
XU_1289 in out fe_tanh Vc=0.3092624635605935 Qo=1.0904318388749068e-13 K=2.62 tau=1.1416994453373934e-07 off=-0.2

*Grain_1290:
XU_1290 in out fe_tanh Vc=0.6601589231192106 Qo=2.3276614310016897e-13 K=2.62 tau=9.888597081994966e-08 off=-0.2

*Grain_1291:
XU_1291 in out fe_tanh Vc=0.23291305483951547 Qo=8.212306393816966e-14 K=2.62 tau=1.0751974087184612e-07 off=-0.2

*Grain_1292:
XU_1292 in out fe_tanh Vc=-0.284465930821407 Qo=1.003001478005343e-13 K=2.62 tau=9.018809496695711e-08 off=-0.2

*Grain_1293:
XU_1293 in out fe_tanh Vc=0.731830971906632 Qo=2.580370676913415e-13 K=2.62 tau=1.0552056020532228e-07 off=-0.2

*Grain_1294:
XU_1294 in out fe_tanh Vc=0.603151972980545 Qo=2.1266600137825716e-13 K=2.62 tau=9.987271432804554e-08 off=-0.2

*Grain_1295:
XU_1295 in out fe_tanh Vc=0.43731406732972106 Qo=1.5419303626894298e-13 K=2.62 tau=1.0428278285425921e-07 off=-0.2

*Grain_1296:
XU_1296 in out fe_tanh Vc=0.6192608903024295 Qo=2.1834586182279657e-13 K=2.62 tau=1.189526998486447e-07 off=-0.2

*Grain_1297:
XU_1297 in out fe_tanh Vc=-0.036194999740662315 Qo=1.2762033798374054e-14 K=2.62 tau=9.914779798208992e-08 off=-0.2

*Grain_1298:
XU_1298 in out fe_tanh Vc=0.3085306232954335 Qo=1.0878514354308116e-13 K=2.62 tau=8.530332505406837e-08 off=-0.2

*Grain_1299:
XU_1299 in out fe_tanh Vc=0.2482848861668782 Qo=8.754303444095488e-14 K=2.62 tau=8.729299327380693e-08 off=-0.2

*Grain_1300:
XU_1300 in out fe_tanh Vc=0.029408136011335684 Qo=1.0369046233262373e-14 K=2.62 tau=1.1265664305047783e-07 off=-0.2

*Grain_1301:
XU_1301 in out fe_tanh Vc=0.6769050405890269 Qo=2.3867067462862884e-13 K=2.62 tau=7.322187154695476e-08 off=-0.2

*Grain_1302:
XU_1302 in out fe_tanh Vc=0.3952068220582924 Qo=1.3934639747461527e-13 K=2.62 tau=9.131778805776817e-08 off=-0.2

*Grain_1303:
XU_1303 in out fe_tanh Vc=0.6329922533737051 Qo=2.2318741786282873e-13 K=2.62 tau=1.2156216706483795e-07 off=-0.2

*Grain_1304:
XU_1304 in out fe_tanh Vc=0.40453920659121695 Qo=1.4263691295139274e-13 K=2.62 tau=1.1159528970646352e-07 off=-0.2

*Grain_1305:
XU_1305 in out fe_tanh Vc=0.3258268639430807 Qo=1.148836435931338e-13 K=2.62 tau=8.948593537928255e-08 off=-0.2

*Grain_1306:
XU_1306 in out fe_tanh Vc=0.41767453418046624 Qo=1.4726831220122869e-13 K=2.62 tau=9.960244596662511e-08 off=-0.2

*Grain_1307:
XU_1307 in out fe_tanh Vc=0.26048138789710534 Qo=9.184341207373113e-14 K=2.62 tau=1.0514695564495389e-07 off=-0.2

*Grain_1308:
XU_1308 in out fe_tanh Vc=0.6441061946250775 Qo=2.2710609433470102e-13 K=2.62 tau=1.1124665789324655e-07 off=-0.2

*Grain_1309:
XU_1309 in out fe_tanh Vc=0.7825012240859912 Qo=2.7590294628005307e-13 K=2.62 tau=9.076686765337156e-08 off=-0.2

*Grain_1310:
XU_1310 in out fe_tanh Vc=0.6274291638198446 Qo=2.2122592214744153e-13 K=2.62 tau=8.781204508313271e-08 off=-0.2

*Grain_1311:
XU_1311 in out fe_tanh Vc=-0.5329725684407942 Qo=1.8792136982408446e-13 K=2.62 tau=9.246279328783883e-08 off=-0.2

*Grain_1312:
XU_1312 in out fe_tanh Vc=0.39082215061562875 Qo=1.378004014655816e-13 K=2.62 tau=1.0739827768853031e-07 off=-0.2

*Grain_1313:
XU_1313 in out fe_tanh Vc=0.7114634553877482 Qo=2.508556631861517e-13 K=2.62 tau=1.033630938175377e-07 off=-0.2

*Grain_1314:
XU_1314 in out fe_tanh Vc=0.19136124452694242 Qo=6.747226655200614e-14 K=2.62 tau=1.2125221974082153e-07 off=-0.2

*Grain_1315:
XU_1315 in out fe_tanh Vc=0.2399725585122924 Qo=8.461218191350457e-14 K=2.62 tau=1.0007660362934489e-07 off=-0.2

*Grain_1316:
XU_1316 in out fe_tanh Vc=0.14940805280031177 Qo=5.267994566234919e-14 K=2.62 tau=8.926660754917281e-08 off=-0.2

*Grain_1317:
XU_1317 in out fe_tanh Vc=0.40843850370924806 Qo=1.4401177030646303e-13 K=2.62 tau=9.248469253853528e-08 off=-0.2

*Grain_1318:
XU_1318 in out fe_tanh Vc=0.58867601672661 Qo=2.075619084289496e-13 K=2.62 tau=9.45221716296742e-08 off=-0.2

*Grain_1319:
XU_1319 in out fe_tanh Vc=0.4839281894517561 Qo=1.7062875960822602e-13 K=2.62 tau=9.954113280646624e-08 off=-0.2

*Grain_1320:
XU_1320 in out fe_tanh Vc=0.43705606702571365 Qo=1.5410206766490032e-13 K=2.62 tau=1.0391047335750164e-07 off=-0.2

*Grain_1321:
XU_1321 in out fe_tanh Vc=0.6615865785013678 Qo=2.3326952164333975e-13 K=2.62 tau=9.817931720555554e-08 off=-0.2

*Grain_1322:
XU_1322 in out fe_tanh Vc=0.1990366035426796 Qo=7.017852962357207e-14 K=2.62 tau=6.777851886582621e-08 off=-0.2

*Grain_1323:
XU_1323 in out fe_tanh Vc=0.3819431556021903 Qo=1.34669747085999e-13 K=2.62 tau=1.1173054503570068e-07 off=-0.2

*Grain_1324:
XU_1324 in out fe_tanh Vc=0.8615267810923858 Qo=3.037666522249916e-13 K=2.62 tau=1.0949318302724541e-07 off=-0.2

*Grain_1325:
XU_1325 in out fe_tanh Vc=0.1502520666881058 Qo=5.2977537424733535e-14 K=2.62 tau=9.635549530788907e-08 off=-0.2

*Grain_1326:
XU_1326 in out fe_tanh Vc=0.5806915604499073 Qo=2.0474666042245645e-13 K=2.62 tau=1.119319378438978e-07 off=-0.2

*Grain_1327:
XU_1327 in out fe_tanh Vc=0.7825290440111903 Qo=2.7591275533733176e-13 K=2.62 tau=8.97917054346136e-08 off=-0.2

*Grain_1328:
XU_1328 in out fe_tanh Vc=0.8551490789317278 Qo=3.0151793137643633e-13 K=2.62 tau=9.887931773645042e-08 off=-0.2

*Grain_1329:
XU_1329 in out fe_tanh Vc=0.25474913727528464 Qo=8.982227167586999e-14 K=2.62 tau=8.926631502036997e-08 off=-0.2

*Grain_1330:
XU_1330 in out fe_tanh Vc=0.08752518458121833 Qo=3.086059875225175e-14 K=2.62 tau=1.027403993942414e-07 off=-0.2

*Grain_1331:
XU_1331 in out fe_tanh Vc=0.5312879235634931 Qo=1.8732737907905284e-13 K=2.62 tau=9.349705034376868e-08 off=-0.2

*Grain_1332:
XU_1332 in out fe_tanh Vc=-0.1390665752213684 Qo=4.9033632985647183e-14 K=2.62 tau=9.73167359382059e-08 off=-0.2

*Grain_1333:
XU_1333 in out fe_tanh Vc=0.0360862960584481 Qo=1.2723705850415345e-14 K=2.62 tau=9.248077758097088e-08 off=-0.2

*Grain_1334:
XU_1334 in out fe_tanh Vc=1.4331017422797037 Qo=5.05298881130691e-13 K=2.62 tau=8.09089898276832e-08 off=-0.2

*Grain_1335:
XU_1335 in out fe_tanh Vc=0.5917295326165325 Qo=2.0863855087321753e-13 K=2.62 tau=8.608647781381509e-08 off=-0.2

*Grain_1336:
XU_1336 in out fe_tanh Vc=0.34087539149090484 Qo=1.2018962006936353e-13 K=2.62 tau=1.05021589906048e-07 off=-0.2

*Grain_1337:
XU_1337 in out fe_tanh Vc=0.4702928760571128 Qo=1.6582106982674582e-13 K=2.62 tau=9.566710563476191e-08 off=-0.2

*Grain_1338:
XU_1338 in out fe_tanh Vc=0.5498001363895746 Qo=1.9385462006432443e-13 K=2.62 tau=7.555382535049095e-08 off=-0.2

*Grain_1339:
XU_1339 in out fe_tanh Vc=0.14323122920474723 Qo=5.050205280261723e-14 K=2.62 tau=1.063467158127544e-07 off=-0.2

*Grain_1340:
XU_1340 in out fe_tanh Vc=0.5063425355142247 Qo=1.7853185793858237e-13 K=2.62 tau=1.0011372570838097e-07 off=-0.2

*Grain_1341:
XU_1341 in out fe_tanh Vc=0.29949833834187467 Qo=1.0560044049902047e-13 K=2.62 tau=1.0075545878934648e-07 off=-0.2

*Grain_1342:
XU_1342 in out fe_tanh Vc=0.36100501045648925 Qo=1.2728714402095448e-13 K=2.62 tau=9.924594197619668e-08 off=-0.2

*Grain_1343:
XU_1343 in out fe_tanh Vc=0.3568103466488471 Qo=1.2580814300784474e-13 K=2.62 tau=1.0239324669237773e-07 off=-0.2

*Grain_1344:
XU_1344 in out fe_tanh Vc=0.42441144902771555 Qo=1.4964368823641e-13 K=2.62 tau=1.0258290307388366e-07 off=-0.2

*Grain_1345:
XU_1345 in out fe_tanh Vc=0.2554307189524896 Qo=9.006259129082138e-14 K=2.62 tau=1.0086810270621829e-07 off=-0.2

*Grain_1346:
XU_1346 in out fe_tanh Vc=0.5439444147514336 Qo=1.9178994488832573e-13 K=2.62 tau=9.120979675494299e-08 off=-0.2

*Grain_1347:
XU_1347 in out fe_tanh Vc=0.936002392098406 Qo=3.3002608782724194e-13 K=2.62 tau=1.1653250162663978e-07 off=-0.2

*Grain_1348:
XU_1348 in out fe_tanh Vc=0.4226937476621394 Qo=1.4903804206870554e-13 K=2.62 tau=1.0004868112010705e-07 off=-0.2

*Grain_1349:
XU_1349 in out fe_tanh Vc=0.464442138154722 Qo=1.6375815187148318e-13 K=2.62 tau=9.679947951379564e-08 off=-0.2

*Grain_1350:
XU_1350 in out fe_tanh Vc=0.39805832631256804 Qo=1.403518124194976e-13 K=2.62 tau=1.0363473998762396e-07 off=-0.2

*Grain_1351:
XU_1351 in out fe_tanh Vc=0.9491052804867695 Qo=3.3464604930442793e-13 K=2.62 tau=1.0662343090759701e-07 off=-0.2

*Grain_1352:
XU_1352 in out fe_tanh Vc=0.2572436438629384 Qo=9.070181243039414e-14 K=2.62 tau=9.644355594487288e-08 off=-0.2

*Grain_1353:
XU_1353 in out fe_tanh Vc=-0.20055358724262456 Qo=7.071340453416728e-14 K=2.62 tau=8.754071185419927e-08 off=-0.2

*Grain_1354:
XU_1354 in out fe_tanh Vc=0.9052605221529468 Qo=3.191867789149554e-13 K=2.62 tau=1.0595906819488511e-07 off=-0.2

*Grain_1355:
XU_1355 in out fe_tanh Vc=-0.08056550365469467 Qo=2.84066773861352e-14 K=2.62 tau=9.631100305581932e-08 off=-0.2

*Grain_1356:
XU_1356 in out fe_tanh Vc=0.13019155590812503 Qo=4.5904380402462564e-14 K=2.62 tau=1.1007461255396286e-07 off=-0.2

*Grain_1357:
XU_1357 in out fe_tanh Vc=0.1889600066263194 Qo=6.66256115039261e-14 K=2.62 tau=9.709180694471451e-08 off=-0.2

*Grain_1358:
XU_1358 in out fe_tanh Vc=-0.06094665801529425 Qo=2.1489247549719623e-14 K=2.62 tau=8.341769466575094e-08 off=-0.2

*Grain_1359:
XU_1359 in out fe_tanh Vc=0.4013052537118101 Qo=1.4149665003538082e-13 K=2.62 tau=9.8867232935475e-08 off=-0.2

*Grain_1360:
XU_1360 in out fe_tanh Vc=0.2460615959065916 Qo=8.675912214233156e-14 K=2.62 tau=9.554509310589423e-08 off=-0.2

*Grain_1361:
XU_1361 in out fe_tanh Vc=0.21079060125507731 Qo=7.432288428986351e-14 K=2.62 tau=9.25119487296862e-08 off=-0.2

*Grain_1362:
XU_1362 in out fe_tanh Vc=0.6508123530243624 Qo=2.294706259208907e-13 K=2.62 tau=9.506730900079488e-08 off=-0.2

*Grain_1363:
XU_1363 in out fe_tanh Vc=0.4890411477230855 Qo=1.7243154305168262e-13 K=2.62 tau=9.83860096433615e-08 off=-0.2

*Grain_1364:
XU_1364 in out fe_tanh Vc=0.18489456340034333 Qo=6.51921725143689e-14 K=2.62 tau=9.568670739027964e-08 off=-0.2

*Grain_1365:
XU_1365 in out fe_tanh Vc=0.027682391195186173 Qo=9.760564016689055e-15 K=2.62 tau=1.0410268257727746e-07 off=-0.2

*Grain_1366:
XU_1366 in out fe_tanh Vc=0.10604220937576214 Qo=3.7389536394647055e-14 K=2.62 tau=9.064132945450443e-08 off=-0.2

*Grain_1367:
XU_1367 in out fe_tanh Vc=0.5086547505670889 Qo=1.7934712432524326e-13 K=2.62 tau=9.072544972119456e-08 off=-0.2

*Grain_1368:
XU_1368 in out fe_tanh Vc=0.4083903298165094 Qo=1.439947846219283e-13 K=2.62 tau=1.0089707726949999e-07 off=-0.2

*Grain_1369:
XU_1369 in out fe_tanh Vc=-0.2871897791167723 Qo=1.0126055239388048e-13 K=2.62 tau=1.066405455335245e-07 off=-0.2

*Grain_1370:
XU_1370 in out fe_tanh Vc=0.46968870337967744 Qo=1.6560804393408855e-13 K=2.62 tau=9.032336542351963e-08 off=-0.2

*Grain_1371:
XU_1371 in out fe_tanh Vc=0.6678700376534862 Qo=2.354850132483846e-13 K=2.62 tau=1.039282279182671e-07 off=-0.2

*Grain_1372:
XU_1372 in out fe_tanh Vc=0.13183905652192224 Qo=4.6485274411766875e-14 K=2.62 tau=1.0494010239665974e-07 off=-0.2

*Grain_1373:
XU_1373 in out fe_tanh Vc=0.14949202198779815 Qo=5.2709552448269934e-14 K=2.62 tau=9.564997835896862e-08 off=-0.2

*Grain_1374:
XU_1374 in out fe_tanh Vc=0.32803773579830425 Qo=1.156631772729901e-13 K=2.62 tau=9.295593517074389e-08 off=-0.2

*Grain_1375:
XU_1375 in out fe_tanh Vc=0.45595669540045364 Qo=1.6076626050527096e-13 K=2.62 tau=1.0046223669945868e-07 off=-0.2

*Grain_1376:
XU_1376 in out fe_tanh Vc=0.6300738571476852 Qo=2.2215841740584923e-13 K=2.62 tau=9.497159894339737e-08 off=-0.2

*Grain_1377:
XU_1377 in out fe_tanh Vc=0.7498157089171342 Qo=2.6437832541277885e-13 K=2.62 tau=9.778606115407137e-08 off=-0.2

*Grain_1378:
XU_1378 in out fe_tanh Vc=0.03174459796786089 Qo=1.1192861861703766e-14 K=2.62 tau=9.371629235648467e-08 off=-0.2

*Grain_1379:
XU_1379 in out fe_tanh Vc=0.18363808831471462 Qo=6.474915061563978e-14 K=2.62 tau=1.132055333756267e-07 off=-0.2

*Grain_1380:
XU_1380 in out fe_tanh Vc=0.4705075521585871 Qo=1.658967627037274e-13 K=2.62 tau=1.0889851344838095e-07 off=-0.2

*Grain_1381:
XU_1381 in out fe_tanh Vc=0.7181337304694214 Qo=2.532075426348793e-13 K=2.62 tau=1.1214898869157886e-07 off=-0.2

*Grain_1382:
XU_1382 in out fe_tanh Vc=0.46905296336901425 Qo=1.6538388768153448e-13 K=2.62 tau=1.0692341495023384e-07 off=-0.2

*Grain_1383:
XU_1383 in out fe_tanh Vc=0.6797243351005235 Qo=2.3966473270574136e-13 K=2.62 tau=9.291215012535448e-08 off=-0.2

*Grain_1384:
XU_1384 in out fe_tanh Vc=0.3811554689456444 Qo=1.3439201580252354e-13 K=2.62 tau=9.962975327544756e-08 off=-0.2

*Grain_1385:
XU_1385 in out fe_tanh Vc=0.6621651837372936 Qo=2.334735326843595e-13 K=2.62 tau=8.401475921436656e-08 off=-0.2

*Grain_1386:
XU_1386 in out fe_tanh Vc=-0.10430709788906506 Qo=3.6777751573654264e-14 K=2.62 tau=9.814758125767906e-08 off=-0.2

*Grain_1387:
XU_1387 in out fe_tanh Vc=0.7039727815700332 Qo=2.482145184667368e-13 K=2.62 tau=9.673385503337388e-08 off=-0.2

*Grain_1388:
XU_1388 in out fe_tanh Vc=0.41506559249205155 Qo=1.4634842265173022e-13 K=2.62 tau=9.380992692822724e-08 off=-0.2

*Grain_1389:
XU_1389 in out fe_tanh Vc=0.2908307012573646 Qo=1.0254430903840083e-13 K=2.62 tau=1.047228413966128e-07 off=-0.2

*Grain_1390:
XU_1390 in out fe_tanh Vc=0.6144928943087923 Qo=2.166647089990006e-13 K=2.62 tau=1.0407126385687656e-07 off=-0.2

*Grain_1391:
XU_1391 in out fe_tanh Vc=0.2837767480590525 Qo=1.0005714811081353e-13 K=2.62 tau=8.671878888006862e-08 off=-0.2

*Grain_1392:
XU_1392 in out fe_tanh Vc=0.57732814918723 Qo=2.0356075163616908e-13 K=2.62 tau=9.379442746267658e-08 off=-0.2

*Grain_1393:
XU_1393 in out fe_tanh Vc=0.2048220127623144 Qo=7.221841326847945e-14 K=2.62 tau=1.2134806349203223e-07 off=-0.2

*Grain_1394:
XU_1394 in out fe_tanh Vc=0.7033583522206508 Qo=2.4799787616311155e-13 K=2.62 tau=8.257789171216216e-08 off=-0.2

*Grain_1395:
XU_1395 in out fe_tanh Vc=0.8950134266483671 Qo=3.15573744515132e-13 K=2.62 tau=1.0889721484778409e-07 off=-0.2

*Grain_1396:
XU_1396 in out fe_tanh Vc=0.03249095616281278 Qo=1.1456021098557381e-14 K=2.62 tau=1.188518881720641e-07 off=-0.2

*Grain_1397:
XU_1397 in out fe_tanh Vc=0.5076516850226824 Qo=1.7899345236858019e-13 K=2.62 tau=9.371023213170686e-08 off=-0.2

*Grain_1398:
XU_1398 in out fe_tanh Vc=0.3751661512277763 Qo=1.3228023584141573e-13 K=2.62 tau=9.388899362522827e-08 off=-0.2

*Grain_1399:
XU_1399 in out fe_tanh Vc=-0.04833285392465092 Qo=1.7041732829889062e-14 K=2.62 tau=9.930709366336247e-08 off=-0.2

*Grain_1400:
XU_1400 in out fe_tanh Vc=-0.19604966430017529 Qo=6.912536151085883e-14 K=2.62 tau=1.0644731077986804e-07 off=-0.2

*Grain_1401:
XU_1401 in out fe_tanh Vc=0.6981940724118013 Qo=2.461769972036691e-13 K=2.62 tau=1.017257530891617e-07 off=-0.2

*Grain_1402:
XU_1402 in out fe_tanh Vc=0.1103526626198661 Qo=3.8909363729409157e-14 K=2.62 tau=1.0596351435398474e-07 off=-0.2

*Grain_1403:
XU_1403 in out fe_tanh Vc=0.6532920495329533 Qo=2.3034494477374585e-13 K=2.62 tau=9.345002109880584e-08 off=-0.2

*Grain_1404:
XU_1404 in out fe_tanh Vc=0.54482781956922 Qo=1.9210142554098533e-13 K=2.62 tau=9.738415813661394e-08 off=-0.2

*Grain_1405:
XU_1405 in out fe_tanh Vc=0.43225700389961713 Qo=1.5240996084753323e-13 K=2.62 tau=9.936314742756392e-08 off=-0.2

*Grain_1406:
XU_1406 in out fe_tanh Vc=0.2725172463666585 Qo=9.608714832684468e-14 K=2.62 tau=9.887719361623094e-08 off=-0.2

*Grain_1407:
XU_1407 in out fe_tanh Vc=0.8772541925997462 Qo=3.093119971250051e-13 K=2.62 tau=1.054485897072966e-07 off=-0.2

*Grain_1408:
XU_1408 in out fe_tanh Vc=0.31666479114367685 Qo=1.1165317851323502e-13 K=2.62 tau=8.951711627662494e-08 off=-0.2

*Grain_1409:
XU_1409 in out fe_tanh Vc=-0.04350863312459924 Qo=1.5340755641266154e-14 K=2.62 tau=9.636761091281159e-08 off=-0.2

*Grain_1410:
XU_1410 in out fe_tanh Vc=0.5196253380120612 Qo=1.8321525552468813e-13 K=2.62 tau=1.0311694351313793e-07 off=-0.2

*Grain_1411:
XU_1411 in out fe_tanh Vc=0.2799615098346472 Qo=9.871192917124797e-14 K=2.62 tau=8.883914265307289e-08 off=-0.2

*Grain_1412:
XU_1412 in out fe_tanh Vc=0.7696454185343073 Qo=2.7137010400538936e-13 K=2.62 tau=1.0995758535884063e-07 off=-0.2

*Grain_1413:
XU_1413 in out fe_tanh Vc=-0.2909817429337049 Qo=1.0259756498514012e-13 K=2.62 tau=9.827748653235006e-08 off=-0.2

*Grain_1414:
XU_1414 in out fe_tanh Vc=0.026853549479304795 Qo=9.468321826680215e-15 K=2.62 tau=9.396822972190163e-08 off=-0.2

*Grain_1415:
XU_1415 in out fe_tanh Vc=0.42575500592629856 Qo=1.5011741440501368e-13 K=2.62 tau=9.194527739401997e-08 off=-0.2

*Grain_1416:
XU_1416 in out fe_tanh Vc=0.35274289340075354 Qo=1.2437399530243228e-13 K=2.62 tau=8.870280037637806e-08 off=-0.2

*Grain_1417:
XU_1417 in out fe_tanh Vc=0.6102270834465534 Qo=2.1516062216956475e-13 K=2.62 tau=1.0617809256852935e-07 off=-0.2

*Grain_1418:
XU_1418 in out fe_tanh Vc=0.1083303458159966 Qo=3.819631287744277e-14 K=2.62 tau=1.0343228125814329e-07 off=-0.2

*Grain_1419:
XU_1419 in out fe_tanh Vc=0.5496363269858427 Qo=1.9379686233088347e-13 K=2.62 tau=9.253356759238322e-08 off=-0.2

*Grain_1420:
XU_1420 in out fe_tanh Vc=0.6473088001751064 Qo=2.2823530446220967e-13 K=2.62 tau=1.1019906424350081e-07 off=-0.2

*Grain_1421:
XU_1421 in out fe_tanh Vc=0.5057984549244341 Qo=1.7834001997959084e-13 K=2.62 tau=8.705658255911991e-08 off=-0.2

*Grain_1422:
XU_1422 in out fe_tanh Vc=0.935056533656458 Qo=3.2969258658422196e-13 K=2.62 tau=8.404885775877068e-08 off=-0.2

*Grain_1423:
XU_1423 in out fe_tanh Vc=0.9184950108807475 Qo=3.238531414970401e-13 K=2.62 tau=8.803032561630815e-08 off=-0.2

*Grain_1424:
XU_1424 in out fe_tanh Vc=0.7753830314946172 Qo=2.733931351159326e-13 K=2.62 tau=1.0825695007547797e-07 off=-0.2

*Grain_1425:
XU_1425 in out fe_tanh Vc=-0.0734142417048827 Qo=2.5885206261437335e-14 K=2.62 tau=9.686636631520794e-08 off=-0.2

*Grain_1426:
XU_1426 in out fe_tanh Vc=0.36113202946868705 Qo=1.2733192979076576e-13 K=2.62 tau=9.134378844831315e-08 off=-0.2

*Grain_1427:
XU_1427 in out fe_tanh Vc=0.4263118750758414 Qo=1.5031376149601127e-13 K=2.62 tau=1.1393225788845915e-07 off=-0.2

*Grain_1428:
XU_1428 in out fe_tanh Vc=0.5237222975706245 Qo=1.8465980689177152e-13 K=2.62 tau=9.703753196715231e-08 off=-0.2

*Grain_1429:
XU_1429 in out fe_tanh Vc=0.3043453679296314 Qo=1.0730945986257574e-13 K=2.62 tau=9.450622023057142e-08 off=-0.2

*Grain_1430:
XU_1430 in out fe_tanh Vc=0.7852258019437586 Qo=2.7686360811058946e-13 K=2.62 tau=9.904473642475478e-08 off=-0.2

*Grain_1431:
XU_1431 in out fe_tanh Vc=0.6556466683218114 Qo=2.3117516233918306e-13 K=2.62 tau=9.971958397528964e-08 off=-0.2

*Grain_1432:
XU_1432 in out fe_tanh Vc=0.17489883382664678 Qo=6.166776749784913e-14 K=2.62 tau=9.77017721247446e-08 off=-0.2

*Grain_1433:
XU_1433 in out fe_tanh Vc=0.8180053043147512 Qo=2.8842136802631953e-13 K=2.62 tau=1.1054482591487546e-07 off=-0.2

*Grain_1434:
XU_1434 in out fe_tanh Vc=0.42174594352005623 Qo=1.4870385478918706e-13 K=2.62 tau=1.1613924641629747e-07 off=-0.2

*Grain_1435:
XU_1435 in out fe_tanh Vc=0.6869359479513886 Qo=2.4220748301940233e-13 K=2.62 tau=1.0852661571198181e-07 off=-0.2

*Grain_1436:
XU_1436 in out fe_tanh Vc=0.39714300169485556 Qo=1.400290771303298e-13 K=2.62 tau=1.0346367457691701e-07 off=-0.2

*Grain_1437:
XU_1437 in out fe_tanh Vc=0.15544902100089986 Qo=5.48099371225839e-14 K=2.62 tau=8.59352077187152e-08 off=-0.2

*Grain_1438:
XU_1438 in out fe_tanh Vc=0.9008491634017541 Qo=3.1763137319917007e-13 K=2.62 tau=8.546957667104381e-08 off=-0.2

*Grain_1439:
XU_1439 in out fe_tanh Vc=0.42000217457968625 Qo=1.4808901742731368e-13 K=2.62 tau=1.0627978794636665e-07 off=-0.2

*Grain_1440:
XU_1440 in out fe_tanh Vc=0.31982904142897617 Qo=1.1276886491679474e-13 K=2.62 tau=1.0646336430454462e-07 off=-0.2

*Grain_1441:
XU_1441 in out fe_tanh Vc=0.9745925745244461 Qo=3.4363264165885503e-13 K=2.62 tau=9.756220923110665e-08 off=-0.2

*Grain_1442:
XU_1442 in out fe_tanh Vc=0.6198714114017566 Qo=2.1856112611234098e-13 K=2.62 tau=8.796735606039982e-08 off=-0.2

*Grain_1443:
XU_1443 in out fe_tanh Vc=0.5161936471291296 Qo=1.8200527195382644e-13 K=2.62 tau=1.1846705004406649e-07 off=-0.2

*Grain_1444:
XU_1444 in out fe_tanh Vc=1.0021177201748785 Qo=3.5333776230018374e-13 K=2.62 tau=1.0197208010727432e-07 off=-0.2

*Grain_1445:
XU_1445 in out fe_tanh Vc=0.24072347415223463 Qo=8.487694806477779e-14 K=2.62 tau=9.517719088678912e-08 off=-0.2

*Grain_1446:
XU_1446 in out fe_tanh Vc=0.1395960871328673 Qo=4.92203341587266e-14 K=2.62 tau=8.50434811839404e-08 off=-0.2

*Grain_1447:
XU_1447 in out fe_tanh Vc=0.19988006988689755 Qo=7.047592832697937e-14 K=2.62 tau=1.1319077028166593e-07 off=-0.2

*Grain_1448:
XU_1448 in out fe_tanh Vc=0.8884234531821604 Qo=3.1325017869917104e-13 K=2.62 tau=9.446296241372177e-08 off=-0.2

*Grain_1449:
XU_1449 in out fe_tanh Vc=0.5347243886071485 Qo=1.885390459763672e-13 K=2.62 tau=9.296568503318393e-08 off=-0.2

*Grain_1450:
XU_1450 in out fe_tanh Vc=0.4069590689433772 Qo=1.434901348148257e-13 K=2.62 tau=1.0769569890183515e-07 off=-0.2

*Grain_1451:
XU_1451 in out fe_tanh Vc=1.0170094289722422 Qo=3.5858844588491085e-13 K=2.62 tau=7.192106045980795e-08 off=-0.2

*Grain_1452:
XU_1452 in out fe_tanh Vc=0.7599779335930985 Qo=2.6796143511606827e-13 K=2.62 tau=8.902529955747629e-08 off=-0.2

*Grain_1453:
XU_1453 in out fe_tanh Vc=0.3474476352194331 Qo=1.2250693453809115e-13 K=2.62 tau=1.1186716862492596e-07 off=-0.2

*Grain_1454:
XU_1454 in out fe_tanh Vc=0.6901511718401298 Qo=2.4334114226049794e-13 K=2.62 tau=1.0652846263589395e-07 off=-0.2

*Grain_1455:
XU_1455 in out fe_tanh Vc=0.23894756036951123 Qo=8.425077671844532e-14 K=2.62 tau=1.1671040878810342e-07 off=-0.2

*Grain_1456:
XU_1456 in out fe_tanh Vc=0.5673337643172667 Qo=2.0003682075018157e-13 K=2.62 tau=1.0380321923942092e-07 off=-0.2

*Grain_1457:
XU_1457 in out fe_tanh Vc=0.29335606736239783 Qo=1.0343473058327228e-13 K=2.62 tau=9.686855603975693e-08 off=-0.2

*Grain_1458:
XU_1458 in out fe_tanh Vc=0.4275983855111554 Qo=1.50767373590916e-13 K=2.62 tau=7.694345768097205e-08 off=-0.2

*Grain_1459:
XU_1459 in out fe_tanh Vc=0.35060485073185754 Qo=1.236201405435341e-13 K=2.62 tau=1.0777962151239694e-07 off=-0.2

*Grain_1460:
XU_1460 in out fe_tanh Vc=0.4611054118280098 Qo=1.625816519554026e-13 K=2.62 tau=8.84411992872721e-08 off=-0.2

*Grain_1461:
XU_1461 in out fe_tanh Vc=0.32540138051160183 Qo=1.1473362193345465e-13 K=2.62 tau=1.003326781733094e-07 off=-0.2

*Grain_1462:
XU_1462 in out fe_tanh Vc=0.5788381598709762 Qo=2.0409316792350023e-13 K=2.62 tau=9.931147487324219e-08 off=-0.2

*Grain_1463:
XU_1463 in out fe_tanh Vc=0.3561951109996003 Qo=1.2559121641008512e-13 K=2.62 tau=1.1581708028214056e-07 off=-0.2

*Grain_1464:
XU_1464 in out fe_tanh Vc=0.24926264601407383 Qo=8.788778383468357e-14 K=2.62 tau=1.0849399317665807e-07 off=-0.2

*Grain_1465:
XU_1465 in out fe_tanh Vc=0.10301093724272326 Qo=3.6320736900487876e-14 K=2.62 tau=1.112716273828808e-07 off=-0.2

*Grain_1466:
XU_1466 in out fe_tanh Vc=0.3255788002239436 Qo=1.147961785402132e-13 K=2.62 tau=9.922812229822725e-08 off=-0.2

*Grain_1467:
XU_1467 in out fe_tanh Vc=0.48569841470416114 Qo=1.7125292522954936e-13 K=2.62 tau=1.0373788974130306e-07 off=-0.2

*Grain_1468:
XU_1468 in out fe_tanh Vc=0.8662063784600857 Qo=3.054166364824104e-13 K=2.62 tau=1.1589585261347661e-07 off=-0.2

*Grain_1469:
XU_1469 in out fe_tanh Vc=0.4074259862494446 Qo=1.436547656888075e-13 K=2.62 tau=1.0104435389412239e-07 off=-0.2

*Grain_1470:
XU_1470 in out fe_tanh Vc=0.15627184197739846 Qo=5.5100056453633084e-14 K=2.62 tau=1.0562677046535729e-07 off=-0.2

*Grain_1471:
XU_1471 in out fe_tanh Vc=0.6468658594251133 Qo=2.2807912750786265e-13 K=2.62 tau=1.0633530919547351e-07 off=-0.2

*Grain_1472:
XU_1472 in out fe_tanh Vc=0.1723093517189614 Qo=6.075473922280152e-14 K=2.62 tau=1.0938407902775332e-07 off=-0.2

*Grain_1473:
XU_1473 in out fe_tanh Vc=0.7496057546736512 Qo=2.643042974207733e-13 K=2.62 tau=1.2052504116628797e-07 off=-0.2

*Grain_1474:
XU_1474 in out fe_tanh Vc=0.5903744306505078 Qo=2.0816075401689588e-13 K=2.62 tau=9.944481906581681e-08 off=-0.2

*Grain_1475:
XU_1475 in out fe_tanh Vc=0.5533705485301358 Qo=1.9511351551227155e-13 K=2.62 tau=1.1903759582484372e-07 off=-0.2

*Grain_1476:
XU_1476 in out fe_tanh Vc=-0.14938216188476588 Qo=5.267081675665407e-14 K=2.62 tau=9.182952245026277e-08 off=-0.2

*Grain_1477:
XU_1477 in out fe_tanh Vc=-0.1187944573254725 Qo=4.188586518330619e-14 K=2.62 tau=9.317318341819871e-08 off=-0.2

*Grain_1478:
XU_1478 in out fe_tanh Vc=0.2783490636622128 Qo=9.814339504503969e-14 K=2.62 tau=1.1471655260676002e-07 off=-0.2

*Grain_1479:
XU_1479 in out fe_tanh Vc=0.05757269289905148 Qo=2.029961756887859e-14 K=2.62 tau=1.1885864495488017e-07 off=-0.2

*Grain_1480:
XU_1480 in out fe_tanh Vc=0.2128870627337451 Qo=7.506207789227954e-14 K=2.62 tau=8.63422365534793e-08 off=-0.2

*Grain_1481:
XU_1481 in out fe_tanh Vc=0.8128594580692521 Qo=2.8660698857675935e-13 K=2.62 tau=1.0791212946144474e-07 off=-0.2

*Grain_1482:
XU_1482 in out fe_tanh Vc=0.45427828028486744 Qo=1.601744663186074e-13 K=2.62 tau=8.71727345981967e-08 off=-0.2

*Grain_1483:
XU_1483 in out fe_tanh Vc=0.7773179078734213 Qo=2.7407535525459534e-13 K=2.62 tau=1.0499062930991651e-07 off=-0.2

*Grain_1484:
XU_1484 in out fe_tanh Vc=0.42196875301651054 Qo=1.4878241542863233e-13 K=2.62 tau=1.0386196764391403e-07 off=-0.2

*Grain_1485:
XU_1485 in out fe_tanh Vc=0.5329953315586301 Qo=1.8792939589622864e-13 K=2.62 tau=1.0927462234187034e-07 off=-0.2

*Grain_1486:
XU_1486 in out fe_tanh Vc=-0.0895592824720855 Qo=3.157780351032459e-14 K=2.62 tau=1.0249304035457076e-07 off=-0.2

*Grain_1487:
XU_1487 in out fe_tanh Vc=0.4866119307584027 Qo=1.715750228353822e-13 K=2.62 tau=1.0613998664691702e-07 off=-0.2

*Grain_1488:
XU_1488 in out fe_tanh Vc=0.5743385705693297 Qo=2.0250665290325274e-13 K=2.62 tau=1.1768205388387438e-07 off=-0.2

*Grain_1489:
XU_1489 in out fe_tanh Vc=0.6923745078539276 Qo=2.441250706914009e-13 K=2.62 tau=9.293769137804222e-08 off=-0.2

*Grain_1490:
XU_1490 in out fe_tanh Vc=0.5188104777239214 Qo=1.8292794306128975e-13 K=2.62 tau=1.0771845189571897e-07 off=-0.2

*Grain_1491:
XU_1491 in out fe_tanh Vc=0.8757925298183203 Qo=3.087966278764338e-13 K=2.62 tau=1.1002319257568418e-07 off=-0.2

*Grain_1492:
XU_1492 in out fe_tanh Vc=1.0527873717348522 Qo=3.712034291158616e-13 K=2.62 tau=9.060592444826678e-08 off=-0.2

*Grain_1493:
XU_1493 in out fe_tanh Vc=0.2861321577862749 Qo=1.0088764455405735e-13 K=2.62 tau=7.970953670523307e-08 off=-0.2

*Grain_1494:
XU_1494 in out fe_tanh Vc=-0.14787311935892172 Qo=5.213874183315651e-14 K=2.62 tau=1.0195337841567094e-07 off=-0.2

*Grain_1495:
XU_1495 in out fe_tanh Vc=0.6640735080419938 Qo=2.341463907987217e-13 K=2.62 tau=9.510251273718195e-08 off=-0.2

*Grain_1496:
XU_1496 in out fe_tanh Vc=1.0493415073559418 Qo=3.6998844809684354e-13 K=2.62 tau=1.024452348768277e-07 off=-0.2

*Grain_1497:
XU_1497 in out fe_tanh Vc=0.40097609497872727 Qo=1.4138059160447236e-13 K=2.62 tau=1.0034610366323293e-07 off=-0.2

*Grain_1498:
XU_1498 in out fe_tanh Vc=0.371655059647864 Qo=1.31042256293603e-13 K=2.62 tau=8.911600383963092e-08 off=-0.2

*Grain_1499:
XU_1499 in out fe_tanh Vc=0.7104379648986917 Qo=2.5049408439419086e-13 K=2.62 tau=9.760897884427508e-08 off=-0.2

*Grain_1500:
XU_1500 in out fe_tanh Vc=0.37315177853885306 Qo=1.3156998601346284e-13 K=2.62 tau=1.1479659328537694e-07 off=-0.2

*Grain_1501:
XU_1501 in out fe_tanh Vc=0.5804981752679976 Qo=2.0467847453365085e-13 K=2.62 tau=1.0766432815787816e-07 off=-0.2

*Grain_1502:
XU_1502 in out fe_tanh Vc=0.48917468050723295 Qo=1.7247862551933536e-13 K=2.62 tau=1.0718955626265982e-07 off=-0.2

*Grain_1503:
XU_1503 in out fe_tanh Vc=0.22806628840127724 Qo=8.041413735878549e-14 K=2.62 tau=1.0083774874727075e-07 off=-0.2

*Grain_1504:
XU_1504 in out fe_tanh Vc=-0.3833151480216082 Qo=1.3515349936540715e-13 K=2.62 tau=9.916073315781025e-08 off=-0.2

*Grain_1505:
XU_1505 in out fe_tanh Vc=0.9225242729774539 Qo=3.252738233434032e-13 K=2.62 tau=1.0291172828126478e-07 off=-0.2

*Grain_1506:
XU_1506 in out fe_tanh Vc=0.12282141575678723 Qo=4.33057347778168e-14 K=2.62 tau=9.272188378892507e-08 off=-0.2

*Grain_1507:
XU_1507 in out fe_tanh Vc=0.5369751175552693 Qo=1.893326329113776e-13 K=2.62 tau=8.791137792738715e-08 off=-0.2

*Grain_1508:
XU_1508 in out fe_tanh Vc=0.6316186961894686 Qo=2.2270311386131402e-13 K=2.62 tau=1.075158976569927e-07 off=-0.2

*Grain_1509:
XU_1509 in out fe_tanh Vc=0.3720476193016417 Qo=1.3118066932317296e-13 K=2.62 tau=1.0756896123946669e-07 off=-0.2

*Grain_1510:
XU_1510 in out fe_tanh Vc=0.8484982553714892 Qo=2.991729103605242e-13 K=2.62 tau=1.1373321041316877e-07 off=-0.2

*Grain_1511:
XU_1511 in out fe_tanh Vc=0.605663953567492 Qo=2.1355170330894298e-13 K=2.62 tau=9.732679569121218e-08 off=-0.2

*Grain_1512:
XU_1512 in out fe_tanh Vc=0.12767292517842516 Qo=4.5016333690807436e-14 K=2.62 tau=1.0148454232847271e-07 off=-0.2

*Grain_1513:
XU_1513 in out fe_tanh Vc=0.6163302848403333 Qo=2.1731255649816756e-13 K=2.62 tau=9.338137822556353e-08 off=-0.2

*Grain_1514:
XU_1514 in out fe_tanh Vc=0.8924433466534023 Qo=3.146675572518283e-13 K=2.62 tau=1.0865475394144906e-07 off=-0.2

*Grain_1515:
XU_1515 in out fe_tanh Vc=0.6198887245859421 Qo=2.1856723058653121e-13 K=2.62 tau=1.2034282374336726e-07 off=-0.2

*Grain_1516:
XU_1516 in out fe_tanh Vc=0.7229107598219509 Qo=2.548918805403806e-13 K=2.62 tau=1.1146346894948443e-07 off=-0.2

*Grain_1517:
XU_1517 in out fe_tanh Vc=0.6105420816321828 Qo=2.1527168771785131e-13 K=2.62 tau=1.2253480302978002e-07 off=-0.2

*Grain_1518:
XU_1518 in out fe_tanh Vc=1.0305870697437955 Qo=3.6337580081432893e-13 K=2.62 tau=1.0307936947283161e-07 off=-0.2

*Grain_1519:
XU_1519 in out fe_tanh Vc=0.45421316470662637 Qo=1.6015150714700173e-13 K=2.62 tau=9.466529582064635e-08 off=-0.2

*Grain_1520:
XU_1520 in out fe_tanh Vc=0.07118777345914218 Qo=2.5100173433512605e-14 K=2.62 tau=7.328460485412062e-08 off=-0.2

*Grain_1521:
XU_1521 in out fe_tanh Vc=0.5387602404701128 Qo=1.8996205131548642e-13 K=2.62 tau=1.012026023993624e-07 off=-0.2

*Grain_1522:
XU_1522 in out fe_tanh Vc=0.024925300521956295 Qo=8.788438457660172e-15 K=2.62 tau=9.326728298978485e-08 off=-0.2

*Grain_1523:
XU_1523 in out fe_tanh Vc=0.41850836453934864 Qo=1.475623133422264e-13 K=2.62 tau=1.0686191003733532e-07 off=-0.2

*Grain_1524:
XU_1524 in out fe_tanh Vc=0.3768922991532553 Qo=1.328888601907401e-13 K=2.62 tau=9.862226017494585e-08 off=-0.2

*Grain_1525:
XU_1525 in out fe_tanh Vc=0.2629500532486961 Qo=9.271384143910235e-14 K=2.62 tau=1.0026507238428104e-07 off=-0.2

*Grain_1526:
XU_1526 in out fe_tanh Vc=0.8632633727698016 Qo=3.043789589480183e-13 K=2.62 tau=8.998848826008063e-08 off=-0.2

*Grain_1527:
XU_1527 in out fe_tanh Vc=0.5505261426102299 Qo=1.9411060337672172e-13 K=2.62 tau=9.315929071824105e-08 off=-0.2

*Grain_1528:
XU_1528 in out fe_tanh Vc=0.5937792723695788 Qo=2.0936127081226093e-13 K=2.62 tau=1.1479926349259997e-07 off=-0.2

*Grain_1529:
XU_1529 in out fe_tanh Vc=0.5180175529706524 Qo=1.826483648716699e-13 K=2.62 tau=1.0239750300080234e-07 off=-0.2

*Grain_1530:
XU_1530 in out fe_tanh Vc=0.2176191314236237 Qo=7.673056306949073e-14 K=2.62 tau=1.00642401504694e-07 off=-0.2

*Grain_1531:
XU_1531 in out fe_tanh Vc=0.8381906559333485 Qo=2.9553854281384146e-13 K=2.62 tau=7.786036536931891e-08 off=-0.2

*Grain_1532:
XU_1532 in out fe_tanh Vc=0.4868254384403387 Qo=1.7165030373806499e-13 K=2.62 tau=1.0757536846008705e-07 off=-0.2

*Grain_1533:
XU_1533 in out fe_tanh Vc=0.6089535733264315 Qo=2.1471159386974387e-13 K=2.62 tau=1.198109285869012e-07 off=-0.2

*Grain_1534:
XU_1534 in out fe_tanh Vc=0.472002003722173 Qo=1.6642369298418517e-13 K=2.62 tau=1.0229936040941826e-07 off=-0.2

*Grain_1535:
XU_1535 in out fe_tanh Vc=0.7721910628594257 Qo=2.7226767546964066e-13 K=2.62 tau=1.0025642885561425e-07 off=-0.2

*Grain_1536:
XU_1536 in out fe_tanh Vc=0.22717653949259078 Qo=8.010041983630775e-14 K=2.62 tau=9.716605612253559e-08 off=-0.2

*Grain_1537:
XU_1537 in out fe_tanh Vc=0.5448549215915263 Qo=1.9211098147211272e-13 K=2.62 tau=9.392666274753585e-08 off=-0.2

*Grain_1538:
XU_1538 in out fe_tanh Vc=0.6089740175682257 Qo=2.1471880232689618e-13 K=2.62 tau=9.625411178791499e-08 off=-0.2

*Grain_1539:
XU_1539 in out fe_tanh Vc=0.1341463837918086 Qo=4.7298817409782686e-14 K=2.62 tau=9.773898105347804e-08 off=-0.2

*Grain_1540:
XU_1540 in out fe_tanh Vc=0.38155944722704305 Qo=1.3453445493825937e-13 K=2.62 tau=1.205642610933997e-07 off=-0.2

*Grain_1541:
XU_1541 in out fe_tanh Vc=0.5901960442441954 Qo=2.0809785656247287e-13 K=2.62 tau=1.0612015980248982e-07 off=-0.2

*Grain_1542:
XU_1542 in out fe_tanh Vc=0.13402689311016258 Qo=4.72566860621191e-14 K=2.62 tau=9.893068095552616e-08 off=-0.2

*Grain_1543:
XU_1543 in out fe_tanh Vc=0.5790929476351312 Qo=2.0418300381466907e-13 K=2.62 tau=9.100228849369279e-08 off=-0.2

*Grain_1544:
XU_1544 in out fe_tanh Vc=0.5617741377493994 Qo=1.980765460527418e-13 K=2.62 tau=1.1494584001490583e-07 off=-0.2

*Grain_1545:
XU_1545 in out fe_tanh Vc=0.41128915356130563 Qo=1.4501688399675043e-13 K=2.62 tau=8.901373727951328e-08 off=-0.2

*Grain_1546:
XU_1546 in out fe_tanh Vc=0.4872370974080832 Qo=1.717954510152414e-13 K=2.62 tau=1.1488780444108627e-07 off=-0.2

*Grain_1547:
XU_1547 in out fe_tanh Vc=1.0626678256409432 Qo=3.746871889610413e-13 K=2.62 tau=7.36539594519216e-08 off=-0.2

*Grain_1548:
XU_1548 in out fe_tanh Vc=0.18230608284789612 Qo=6.427949737875748e-14 K=2.62 tau=1.0403758676974567e-07 off=-0.2

*Grain_1549:
XU_1549 in out fe_tanh Vc=0.9059745777386607 Qo=3.194385485401548e-13 K=2.62 tau=1.05591040689584e-07 off=-0.2

*Grain_1550:
XU_1550 in out fe_tanh Vc=0.07542996104778898 Qo=2.6595930907563155e-14 K=2.62 tau=9.954850198468012e-08 off=-0.2

*Grain_1551:
XU_1551 in out fe_tanh Vc=0.38355842814995983 Qo=1.3523927776691958e-13 K=2.62 tau=1.083071862493132e-07 off=-0.2

*Grain_1552:
XU_1552 in out fe_tanh Vc=0.27331567503901355 Qo=9.63686671492012e-14 K=2.62 tau=9.750897452196378e-08 off=-0.2

*Grain_1553:
XU_1553 in out fe_tanh Vc=0.09866670396310506 Qo=3.4788999026755416e-14 K=2.62 tau=9.677950640457661e-08 off=-0.2

*Grain_1554:
XU_1554 in out fe_tanh Vc=0.38587326606842287 Qo=1.360554689525765e-13 K=2.62 tau=1.0314135350137145e-07 off=-0.2

*Grain_1555:
XU_1555 in out fe_tanh Vc=0.9906562939487178 Qo=3.492965657281746e-13 K=2.62 tau=1.112607602375317e-07 off=-0.2

*Grain_1556:
XU_1556 in out fe_tanh Vc=0.4041898667542706 Qo=1.4251373884341733e-13 K=2.62 tau=1.1618916541931418e-07 off=-0.2

*Grain_1557:
XU_1557 in out fe_tanh Vc=0.8550023816635905 Qo=3.0146620722924715e-13 K=2.62 tau=1.210308275153196e-07 off=-0.2

*Grain_1558:
XU_1558 in out fe_tanh Vc=0.48620531654918786 Qo=1.714316542950291e-13 K=2.62 tau=9.861537584633831e-08 off=-0.2

*Grain_1559:
XU_1559 in out fe_tanh Vc=0.1487759974025606 Qo=5.2457088571415624e-14 K=2.62 tau=9.714665002009004e-08 off=-0.2

*Grain_1560:
XU_1560 in out fe_tanh Vc=0.39555816308085634 Qo=1.3947027718277506e-13 K=2.62 tau=8.611557424182706e-08 off=-0.2

*Grain_1561:
XU_1561 in out fe_tanh Vc=0.2675156114734516 Qo=9.432361651273821e-14 K=2.62 tau=1.127264933110889e-07 off=-0.2

*Grain_1562:
XU_1562 in out fe_tanh Vc=0.3102191561911734 Qo=1.0938050516870621e-13 K=2.62 tau=7.99169184104843e-08 off=-0.2

*Grain_1563:
XU_1563 in out fe_tanh Vc=0.30533676036792534 Qo=1.0765901598622854e-13 K=2.62 tau=8.979902123114188e-08 off=-0.2

*Grain_1564:
XU_1564 in out fe_tanh Vc=0.378019383230729 Qo=1.3328625997505808e-13 K=2.62 tau=1.0984714042209157e-07 off=-0.2

*Grain_1565:
XU_1565 in out fe_tanh Vc=0.15058159910399832 Qo=5.309372761286484e-14 K=2.62 tau=9.604236291831131e-08 off=-0.2

*Grain_1566:
XU_1566 in out fe_tanh Vc=1.0711173031344654 Qo=3.776663992973737e-13 K=2.62 tau=1.1129760068686951e-07 off=-0.2

*Grain_1567:
XU_1567 in out fe_tanh Vc=0.038413779136923176 Qo=1.354435560661007e-14 K=2.62 tau=9.542201778718128e-08 off=-0.2

*Grain_1568:
XU_1568 in out fe_tanh Vc=0.5355699038002242 Qo=1.8883716708559178e-13 K=2.62 tau=9.18311362171871e-08 off=-0.2

*Grain_1569:
XU_1569 in out fe_tanh Vc=-0.5011653457731664 Qo=1.7670642705228911e-13 K=2.62 tau=9.204942653089942e-08 off=-0.2

*Grain_1570:
XU_1570 in out fe_tanh Vc=0.8058156200694597 Qo=2.8412339417787245e-13 K=2.62 tau=1.0689222553640068e-07 off=-0.2

*Grain_1571:
XU_1571 in out fe_tanh Vc=0.563208860006128 Qo=1.9858241631280096e-13 K=2.62 tau=9.589548373001302e-08 off=-0.2

*Grain_1572:
XU_1572 in out fe_tanh Vc=0.538643468028583 Qo=1.8992087839502226e-13 K=2.62 tau=8.921291245644633e-08 off=-0.2

*Grain_1573:
XU_1573 in out fe_tanh Vc=0.6774473032770187 Qo=2.388618716116744e-13 K=2.62 tau=9.984440819611059e-08 off=-0.2

*Grain_1574:
XU_1574 in out fe_tanh Vc=0.2816708498136878 Qo=9.93146271887015e-14 K=2.62 tau=1.1044839475522515e-07 off=-0.2

*Grain_1575:
XU_1575 in out fe_tanh Vc=0.48391226921869007 Qo=1.7062314627616572e-13 K=2.62 tau=1.2093620931270115e-07 off=-0.2

*Grain_1576:
XU_1576 in out fe_tanh Vc=1.3536960905527147 Qo=4.773011571803493e-13 K=2.62 tau=9.413397011950252e-08 off=-0.2

*Grain_1577:
XU_1577 in out fe_tanh Vc=0.711785082612785 Qo=2.509690660745563e-13 K=2.62 tau=9.1057959247585e-08 off=-0.2

*Grain_1578:
XU_1578 in out fe_tanh Vc=0.5561353996903277 Qo=1.9608837734972593e-13 K=2.62 tau=9.553144185349238e-08 off=-0.2

*Grain_1579:
XU_1579 in out fe_tanh Vc=0.6301728408666569 Qo=2.2219331818153805e-13 K=2.62 tau=9.01073579480424e-08 off=-0.2

*Grain_1580:
XU_1580 in out fe_tanh Vc=-0.018323808630545613 Qo=6.460811347796468e-15 K=2.62 tau=1.1239559355094332e-07 off=-0.2

*Grain_1581:
XU_1581 in out fe_tanh Vc=0.24733636871058798 Qo=8.720859565321469e-14 K=2.62 tau=9.43113407248268e-08 off=-0.2

*Grain_1582:
XU_1582 in out fe_tanh Vc=0.4914247168540181 Qo=1.732719682492977e-13 K=2.62 tau=1.2307226219187607e-07 off=-0.2

*Grain_1583:
XU_1583 in out fe_tanh Vc=0.5325924745284112 Qo=1.8778735210364948e-13 K=2.62 tau=1.1324534553750947e-07 off=-0.2

*Grain_1584:
XU_1584 in out fe_tanh Vc=-0.041557272327200634 Qo=1.4652723243762193e-14 K=2.62 tau=1.0390061700926974e-07 off=-0.2

*Grain_1585:
XU_1585 in out fe_tanh Vc=0.47856472841978337 Qo=1.6873765112758688e-13 K=2.62 tau=1.0884211998667911e-07 off=-0.2

*Grain_1586:
XU_1586 in out fe_tanh Vc=0.5176942166076669 Qo=1.8253435935648186e-13 K=2.62 tau=9.15864223542871e-08 off=-0.2

*Grain_1587:
XU_1587 in out fe_tanh Vc=0.7774244648278892 Qo=2.741129262855144e-13 K=2.62 tau=9.990260316088595e-08 off=-0.2

*Grain_1588:
XU_1588 in out fe_tanh Vc=0.49207640988886114 Qo=1.7350174939576604e-13 K=2.62 tau=6.863786406360891e-08 off=-0.2

*Grain_1589:
XU_1589 in out fe_tanh Vc=0.4732056207769522 Qo=1.6684807761309664e-13 K=2.62 tau=1.0523436314109506e-07 off=-0.2

*Grain_1590:
XU_1590 in out fe_tanh Vc=0.15677154858684827 Qo=5.527624854327979e-14 K=2.62 tau=1.1495071071762475e-07 off=-0.2

*Grain_1591:
XU_1591 in out fe_tanh Vc=0.43347433267975066 Qo=1.5283918010840103e-13 K=2.62 tau=9.976702573582939e-08 off=-0.2

*Grain_1592:
XU_1592 in out fe_tanh Vc=0.5389382052539433 Qo=1.900248001095861e-13 K=2.62 tau=8.771538906379025e-08 off=-0.2

*Grain_1593:
XU_1593 in out fe_tanh Vc=0.04904491204746925 Qo=1.7292798167502682e-14 K=2.62 tau=9.518770545680147e-08 off=-0.2

*Grain_1594:
XU_1594 in out fe_tanh Vc=0.3950059763381776 Qo=1.3927558106663822e-13 K=2.62 tau=1.0102933204592583e-07 off=-0.2

*Grain_1595:
XU_1595 in out fe_tanh Vc=0.7578404952672906 Qo=2.6720779344314807e-13 K=2.62 tau=1.0952885857455142e-07 off=-0.2

*Grain_1596:
XU_1596 in out fe_tanh Vc=0.29935949553165775 Qo=1.0555148576357786e-13 K=2.62 tau=8.291249074400028e-08 off=-0.2

*Grain_1597:
XU_1597 in out fe_tanh Vc=0.18425278552722685 Qo=6.496588736541339e-14 K=2.62 tau=1.073073038108855e-07 off=-0.2

*Grain_1598:
XU_1598 in out fe_tanh Vc=0.2767227064188449 Qo=9.756995599940338e-14 K=2.62 tau=9.352029931244529e-08 off=-0.2

*Grain_1599:
XU_1599 in out fe_tanh Vc=0.6622605647486226 Qo=2.335071631774946e-13 K=2.62 tau=1.0784567125696262e-07 off=-0.2

*Grain_1600:
XU_1600 in out fe_tanh Vc=-0.27002176898004465 Qo=9.520726527727344e-14 K=2.62 tau=9.53556373946572e-08 off=-0.2

*Grain_1601:
XU_1601 in out fe_tanh Vc=0.5531734483290466 Qo=1.9504401974086697e-13 K=2.62 tau=9.194239084863916e-08 off=-0.2

*Grain_1602:
XU_1602 in out fe_tanh Vc=0.7916916224422951 Qo=2.7914339869845453e-13 K=2.62 tau=9.969807968613276e-08 off=-0.2

*Grain_1603:
XU_1603 in out fe_tanh Vc=0.10560204453728578 Qo=3.723433820192043e-14 K=2.62 tau=1.1758781265790496e-07 off=-0.2

*Grain_1604:
XU_1604 in out fe_tanh Vc=0.8506744507527908 Qo=2.9994021742523e-13 K=2.62 tau=1.0664575803426006e-07 off=-0.2

*Grain_1605:
XU_1605 in out fe_tanh Vc=0.2794298609061947 Qo=9.852447450506772e-14 K=2.62 tau=9.498173558458916e-08 off=-0.2

*Grain_1606:
XU_1606 in out fe_tanh Vc=0.6401092086334996 Qo=2.256967927548798e-13 K=2.62 tau=1.1110749980513785e-07 off=-0.2

*Grain_1607:
XU_1607 in out fe_tanh Vc=0.0920042351232373 Qo=3.2439871989202624e-14 K=2.62 tau=1.121296226874737e-07 off=-0.2

*Grain_1608:
XU_1608 in out fe_tanh Vc=0.2857311872544709 Qo=1.0074626592397863e-13 K=2.62 tau=8.529179084428816e-08 off=-0.2

*Grain_1609:
XU_1609 in out fe_tanh Vc=0.5951550671252621 Qo=2.098463637614931e-13 K=2.62 tau=1.1953089058300916e-07 off=-0.2

*Grain_1610:
XU_1610 in out fe_tanh Vc=0.3333970297712607 Qo=1.1755281648581915e-13 K=2.62 tau=1.0581124504544443e-07 off=-0.2

*Grain_1611:
XU_1611 in out fe_tanh Vc=0.9871811842696039 Qo=3.4807127307737556e-13 K=2.62 tau=9.623609860862541e-08 off=-0.2

*Grain_1612:
XU_1612 in out fe_tanh Vc=0.5906705512367845 Qo=2.0826516349216966e-13 K=2.62 tau=9.475940212067306e-08 off=-0.2

*Grain_1613:
XU_1613 in out fe_tanh Vc=0.8378746287835132 Qo=2.954271144619614e-13 K=2.62 tau=1.0916522371473138e-07 off=-0.2

*Grain_1614:
XU_1614 in out fe_tanh Vc=0.44866138255450894 Qo=1.5819399832052878e-13 K=2.62 tau=1.1921473663063963e-07 off=-0.2

*Grain_1615:
XU_1615 in out fe_tanh Vc=0.7243966516717053 Qo=2.554157927421533e-13 K=2.62 tau=8.989456209084738e-08 off=-0.2

*Grain_1616:
XU_1616 in out fe_tanh Vc=0.11461646732604402 Qo=4.0412743206126716e-14 K=2.62 tau=9.576585976506475e-08 off=-0.2

*Grain_1617:
XU_1617 in out fe_tanh Vc=0.2558294230431529 Qo=9.020317079398626e-14 K=2.62 tau=1.0835905269922518e-07 off=-0.2

*Grain_1618:
XU_1618 in out fe_tanh Vc=0.5794352043411033 Qo=2.0430368047389363e-13 K=2.62 tau=9.039056226553945e-08 off=-0.2

*Grain_1619:
XU_1619 in out fe_tanh Vc=0.7462417411089035 Qo=2.631181762681527e-13 K=2.62 tau=8.797736647257464e-08 off=-0.2

*Grain_1620:
XU_1620 in out fe_tanh Vc=0.39346562614780334 Qo=1.3873246734010863e-13 K=2.62 tau=1.0771542400987845e-07 off=-0.2

*Grain_1621:
XU_1621 in out fe_tanh Vc=0.6910776940298887 Qo=2.436678257136094e-13 K=2.62 tau=9.363151506945964e-08 off=-0.2

*Grain_1622:
XU_1622 in out fe_tanh Vc=0.7802731232083535 Qo=2.7511733780069577e-13 K=2.62 tau=9.795658813587578e-08 off=-0.2

*Grain_1623:
XU_1623 in out fe_tanh Vc=0.7936850405474462 Qo=2.798462601272294e-13 K=2.62 tau=1.0145457406433789e-07 off=-0.2

*Grain_1624:
XU_1624 in out fe_tanh Vc=0.384496403331821 Qo=1.3556999944280623e-13 K=2.62 tau=9.816175418644661e-08 off=-0.2

*Grain_1625:
XU_1625 in out fe_tanh Vc=0.8533141381127801 Qo=3.008709476240613e-13 K=2.62 tau=1.1066555327140676e-07 off=-0.2

*Grain_1626:
XU_1626 in out fe_tanh Vc=0.3814438602472695 Qo=1.3449370000102797e-13 K=2.62 tau=9.723619562020302e-08 off=-0.2

*Grain_1627:
XU_1627 in out fe_tanh Vc=0.05495354929591667 Qo=1.937613091532157e-14 K=2.62 tau=8.254325265630675e-08 off=-0.2

*Grain_1628:
XU_1628 in out fe_tanh Vc=0.6129292394394003 Qo=2.1611337825068852e-13 K=2.62 tau=9.422265265204617e-08 off=-0.2

*Grain_1629:
XU_1629 in out fe_tanh Vc=0.7330897350180365 Qo=2.5848089632753415e-13 K=2.62 tau=1.0474545054312371e-07 off=-0.2

*Grain_1630:
XU_1630 in out fe_tanh Vc=0.37600868473893034 Qo=1.3257730563621205e-13 K=2.62 tau=9.646055151374942e-08 off=-0.2

*Grain_1631:
XU_1631 in out fe_tanh Vc=0.031719739478961395 Qo=1.1184096980427763e-14 K=2.62 tau=1.0381282016714149e-07 off=-0.2

*Grain_1632:
XU_1632 in out fe_tanh Vc=0.46246023106082 Qo=1.6305934912251674e-13 K=2.62 tau=8.879506427402371e-08 off=-0.2

*Grain_1633:
XU_1633 in out fe_tanh Vc=0.9207410102462239 Qo=3.2464506082343083e-13 K=2.62 tau=1.2356185781115109e-07 off=-0.2

*Grain_1634:
XU_1634 in out fe_tanh Vc=0.4577104529584905 Qo=1.61384619764566e-13 K=2.62 tau=9.746048015305698e-08 off=-0.2

*Grain_1635:
XU_1635 in out fe_tanh Vc=0.2896511795700733 Qo=1.0212842022096796e-13 K=2.62 tau=9.19986546225569e-08 off=-0.2

*Grain_1636:
XU_1636 in out fe_tanh Vc=0.34375927610933255 Qo=1.2120645204158862e-13 K=2.62 tau=9.063707323560107e-08 off=-0.2

*Grain_1637:
XU_1637 in out fe_tanh Vc=1.3005627598840335 Qo=4.58566819104029e-13 K=2.62 tau=1.0424569822583272e-07 off=-0.2

*Grain_1638:
XU_1638 in out fe_tanh Vc=0.722595824162221 Qo=2.54780837038168e-13 K=2.62 tau=8.14121747359319e-08 off=-0.2

*Grain_1639:
XU_1639 in out fe_tanh Vc=0.2843884282860165 Qo=1.0027282109841523e-13 K=2.62 tau=9.988170149241513e-08 off=-0.2

*Grain_1640:
XU_1640 in out fe_tanh Vc=0.2822793312967167 Qo=9.952917232774664e-14 K=2.62 tau=1.1279193254449491e-07 off=-0.2

*Grain_1641:
XU_1641 in out fe_tanh Vc=0.6450286186984191 Qo=2.274313328285473e-13 K=2.62 tau=9.510729112803122e-08 off=-0.2

*Grain_1642:
XU_1642 in out fe_tanh Vc=0.46558522857598766 Qo=1.641611953497347e-13 K=2.62 tau=1.1032383150203558e-07 off=-0.2

*Grain_1643:
XU_1643 in out fe_tanh Vc=1.035887387103303 Qo=3.6524464539973587e-13 K=2.62 tau=9.689631376583376e-08 off=-0.2

*Grain_1644:
XU_1644 in out fe_tanh Vc=0.250222024789962 Qo=8.822605222675578e-14 K=2.62 tau=9.328726507067472e-08 off=-0.2

*Grain_1645:
XU_1645 in out fe_tanh Vc=0.5030257723124189 Qo=1.7736239684213437e-13 K=2.62 tau=1.0659075296108612e-07 off=-0.2

*Grain_1646:
XU_1646 in out fe_tanh Vc=0.18872389452257748 Qo=6.654236048390263e-14 K=2.62 tau=1.0617888854455438e-07 off=-0.2

*Grain_1647:
XU_1647 in out fe_tanh Vc=1.1903115433225575 Qo=4.196932243492065e-13 K=2.62 tau=1.0317852661063803e-07 off=-0.2

*Grain_1648:
XU_1648 in out fe_tanh Vc=0.7233592468251133 Qo=2.5505001305408415e-13 K=2.62 tau=8.839051072247728e-08 off=-0.2

*Grain_1649:
XU_1649 in out fe_tanh Vc=0.09990077680737897 Qo=3.522412209516605e-14 K=2.62 tau=9.245034659559678e-08 off=-0.2

*Grain_1650:
XU_1650 in out fe_tanh Vc=-0.11834590554195296 Qo=4.1727709828627003e-14 K=2.62 tau=8.863607172507935e-08 off=-0.2

*Grain_1651:
XU_1651 in out fe_tanh Vc=0.030313589540985786 Qo=1.068830106489786e-14 K=2.62 tau=8.431942239928801e-08 off=-0.2

*Grain_1652:
XU_1652 in out fe_tanh Vc=0.8891644634576434 Qo=3.135114523073604e-13 K=2.62 tau=1.037076981148181e-07 off=-0.2

*Grain_1653:
XU_1653 in out fe_tanh Vc=0.6908672544992465 Qo=2.435936266136836e-13 K=2.62 tau=9.702685229589826e-08 off=-0.2

*Grain_1654:
XU_1654 in out fe_tanh Vc=0.618492629998653 Qo=2.1807498009788995e-13 K=2.62 tau=1.1123508104310305e-07 off=-0.2

*Grain_1655:
XU_1655 in out fe_tanh Vc=0.38017283216970266 Qo=1.3404554684725497e-13 K=2.62 tau=7.64046761157341e-08 off=-0.2

*Grain_1656:
XU_1656 in out fe_tanh Vc=0.4061284549157861 Qo=1.431972677235293e-13 K=2.62 tau=9.98997160154813e-08 off=-0.2

*Grain_1657:
XU_1657 in out fe_tanh Vc=1.1095711213180335 Qo=3.9122487231440507e-13 K=2.62 tau=9.813447474438515e-08 off=-0.2

*Grain_1658:
XU_1658 in out fe_tanh Vc=1.362701574061313 Qo=4.804764102741716e-13 K=2.62 tau=9.808069088492219e-08 off=-0.2

*Grain_1659:
XU_1659 in out fe_tanh Vc=1.0775939553512337 Qo=3.799500090523934e-13 K=2.62 tau=9.232158138404241e-08 off=-0.2

*Grain_1660:
XU_1660 in out fe_tanh Vc=0.09293520581419423 Qo=3.276812394412501e-14 K=2.62 tau=9.308201460737662e-08 off=-0.2

*Grain_1661:
XU_1661 in out fe_tanh Vc=0.968192472912569 Qo=3.4137602296375824e-13 K=2.62 tau=1.0462158917336238e-07 off=-0.2

*Grain_1662:
XU_1662 in out fe_tanh Vc=0.017320710820041885 Qo=6.107128014395527e-15 K=2.62 tau=8.427698683078787e-08 off=-0.2

*Grain_1663:
XU_1663 in out fe_tanh Vc=0.7428423300553704 Qo=2.619195742769771e-13 K=2.62 tau=9.682901506026658e-08 off=-0.2

*Grain_1664:
XU_1664 in out fe_tanh Vc=0.12573803378697762 Qo=4.433410825882061e-14 K=2.62 tau=8.66560366754055e-08 off=-0.2

*Grain_1665:
XU_1665 in out fe_tanh Vc=0.05828763543612164 Qo=2.055169992520845e-14 K=2.62 tau=9.491442746590919e-08 off=-0.2

*Grain_1666:
XU_1666 in out fe_tanh Vc=0.7211709345818702 Qo=2.542784336920241e-13 K=2.62 tau=1.0125463602866957e-07 off=-0.2

*Grain_1667:
XU_1667 in out fe_tanh Vc=0.8203779901309582 Qo=2.89257955864317e-13 K=2.62 tau=1.2190699812237596e-07 off=-0.2

*Grain_1668:
XU_1668 in out fe_tanh Vc=0.06825899870423013 Qo=2.4067513599894152e-14 K=2.62 tau=1.0556364462140368e-07 off=-0.2

*Grain_1669:
XU_1669 in out fe_tanh Vc=1.3899326475507292 Qo=4.900778436966871e-13 K=2.62 tau=9.432743230236693e-08 off=-0.2

*Grain_1670:
XU_1670 in out fe_tanh Vc=0.4331021448303328 Qo=1.5270794999519072e-13 K=2.62 tau=1.2115041135801034e-07 off=-0.2

*Grain_1671:
XU_1671 in out fe_tanh Vc=0.8034985366325129 Qo=2.8330641124244377e-13 K=2.62 tau=9.717867464114163e-08 off=-0.2

*Grain_1672:
XU_1672 in out fe_tanh Vc=0.04459444566030357 Qo=1.572360344838437e-14 K=2.62 tau=8.916099373378536e-08 off=-0.2

*Grain_1673:
XU_1673 in out fe_tanh Vc=1.0206734280147565 Qo=3.59880339239043e-13 K=2.62 tau=9.926377014122659e-08 off=-0.2

*Grain_1674:
XU_1674 in out fe_tanh Vc=0.21998695180095162 Qo=7.756543539717277e-14 K=2.62 tau=8.503452558059716e-08 off=-0.2

*Grain_1675:
XU_1675 in out fe_tanh Vc=0.5105841252582567 Qo=1.8002740461795865e-13 K=2.62 tau=9.823041165216194e-08 off=-0.2

*Grain_1676:
XU_1676 in out fe_tanh Vc=0.36394519303653705 Qo=1.2832382615187896e-13 K=2.62 tau=8.834306724770302e-08 off=-0.2

*Grain_1677:
XU_1677 in out fe_tanh Vc=0.5933909173246508 Qo=2.0922434029023712e-13 K=2.62 tau=9.363928537628451e-08 off=-0.2

*Grain_1678:
XU_1678 in out fe_tanh Vc=0.6809936994198066 Qo=2.4011229923319574e-13 K=2.62 tau=9.846260676549242e-08 off=-0.2

*Grain_1679:
XU_1679 in out fe_tanh Vc=0.3250325520804131 Qo=1.146035763211226e-13 K=2.62 tau=1.0757613858660296e-07 off=-0.2

*Grain_1680:
XU_1680 in out fe_tanh Vc=0.4183748653359403 Qo=1.475152427148425e-13 K=2.62 tau=9.404344528642666e-08 off=-0.2

*Grain_1681:
XU_1681 in out fe_tanh Vc=0.2996966661323138 Qo=1.0567036910747126e-13 K=2.62 tau=1.0354234507749275e-07 off=-0.2

*Grain_1682:
XU_1682 in out fe_tanh Vc=0.14166149553450835 Qo=4.9948578723391605e-14 K=2.62 tau=9.866652654643351e-08 off=-0.2

*Grain_1683:
XU_1683 in out fe_tanh Vc=0.7421714739334079 Qo=2.616830363970579e-13 K=2.62 tau=1.0579818088028973e-07 off=-0.2

*Grain_1684:
XU_1684 in out fe_tanh Vc=1.0280246934475135 Qo=3.6247232980641045e-13 K=2.62 tau=1.0694187474752764e-07 off=-0.2

*Grain_1685:
XU_1685 in out fe_tanh Vc=0.21288553502883853 Qo=7.506153923716719e-14 K=2.62 tau=1.1402323018710192e-07 off=-0.2

*Grain_1686:
XU_1686 in out fe_tanh Vc=0.48371999359341566 Qo=1.705553516071248e-13 K=2.62 tau=9.736289084072987e-08 off=-0.2

*Grain_1687:
XU_1687 in out fe_tanh Vc=0.44822415506668395 Qo=1.5803983581142032e-13 K=2.62 tau=1.0159009439289161e-07 off=-0.2

*Grain_1688:
XU_1688 in out fe_tanh Vc=0.24131279739763875 Qo=8.508473818026067e-14 K=2.62 tau=8.77491857569827e-08 off=-0.2

*Grain_1689:
XU_1689 in out fe_tanh Vc=0.7950765945957277 Qo=2.8033690966234967e-13 K=2.62 tau=9.829423753743917e-08 off=-0.2

*Grain_1690:
XU_1690 in out fe_tanh Vc=0.3633048751326975 Qo=1.2809805577505744e-13 K=2.62 tau=1.2095480924514347e-07 off=-0.2

*Grain_1691:
XU_1691 in out fe_tanh Vc=0.9710945831839974 Qo=3.4239928113853224e-13 K=2.62 tau=9.582961713294021e-08 off=-0.2

*Grain_1692:
XU_1692 in out fe_tanh Vc=0.3141673323180238 Qo=1.1077259682594671e-13 K=2.62 tau=9.070197986477142e-08 off=-0.2

*Grain_1693:
XU_1693 in out fe_tanh Vc=0.3310974727335148 Qo=1.1674201320229178e-13 K=2.62 tau=1.2146475897992313e-07 off=-0.2

*Grain_1694:
XU_1694 in out fe_tanh Vc=0.049834430894705795 Qo=1.7571175465059796e-14 K=2.62 tau=1.0269729351541239e-07 off=-0.2

*Grain_1695:
XU_1695 in out fe_tanh Vc=0.5537025529444685 Qo=1.9523057730498552e-13 K=2.62 tau=9.836162447540515e-08 off=-0.2

*Grain_1696:
XU_1696 in out fe_tanh Vc=0.26357338783260775 Qo=9.293362364892619e-14 K=2.62 tau=1.0042992939448401e-07 off=-0.2

*Grain_1697:
XU_1697 in out fe_tanh Vc=0.8551676473833774 Qo=3.015244784467287e-13 K=2.62 tau=1.1080132464577056e-07 off=-0.2

*Grain_1698:
XU_1698 in out fe_tanh Vc=0.5054097128384323 Qo=1.782029529903395e-13 K=2.62 tau=1.0292664269102633e-07 off=-0.2

*Grain_1699:
XU_1699 in out fe_tanh Vc=0.6744800950415787 Qo=2.378156604759147e-13 K=2.62 tau=9.679331773789034e-08 off=-0.2

*Grain_1700:
XU_1700 in out fe_tanh Vc=0.17866521257376278 Qo=6.299575902188754e-14 K=2.62 tau=1.0407716616497325e-07 off=-0.2

*Grain_1701:
XU_1701 in out fe_tanh Vc=0.2560949761796172 Qo=9.029680245932963e-14 K=2.62 tau=9.059325577094637e-08 off=-0.2

*Grain_1702:
XU_1702 in out fe_tanh Vc=0.5998193464058013 Qo=2.1149094699812244e-13 K=2.62 tau=1.1045578795957865e-07 off=-0.2

*Grain_1703:
XU_1703 in out fe_tanh Vc=0.41973338215097816 Qo=1.4799424361644207e-13 K=2.62 tau=9.748108962159778e-08 off=-0.2

*Grain_1704:
XU_1704 in out fe_tanh Vc=0.2449046709557713 Qo=8.63512007324589e-14 K=2.62 tau=8.560565095574969e-08 off=-0.2

*Grain_1705:
XU_1705 in out fe_tanh Vc=0.5972541093773527 Qo=2.1058646732157964e-13 K=2.62 tau=9.475439801743166e-08 off=-0.2

*Grain_1706:
XU_1706 in out fe_tanh Vc=-0.19824088126817813 Qo=6.98979650529389e-14 K=2.62 tau=8.917260559984802e-08 off=-0.2

*Grain_1707:
XU_1707 in out fe_tanh Vc=-0.03615139655666272 Qo=1.2746659704938311e-14 K=2.62 tau=1.1958910988642482e-07 off=-0.2

*Grain_1708:
XU_1708 in out fe_tanh Vc=0.7247728393722824 Qo=2.55548433167176e-13 K=2.62 tau=9.792431805178123e-08 off=-0.2

*Grain_1709:
XU_1709 in out fe_tanh Vc=-0.17431777597823678 Qo=6.146289168756178e-14 K=2.62 tau=1.0253887941291654e-07 off=-0.2

*Grain_1710:
XU_1710 in out fe_tanh Vc=0.5780284398082725 Qo=2.0380766785770422e-13 K=2.62 tau=9.72469256966049e-08 off=-0.2

*Grain_1711:
XU_1711 in out fe_tanh Vc=0.7111457860771007 Qo=2.5074365582302863e-13 K=2.62 tau=8.084982640107578e-08 off=-0.2

*Grain_1712:
XU_1712 in out fe_tanh Vc=0.3323433597058371 Qo=1.171813018267884e-13 K=2.62 tau=9.039252781269731e-08 off=-0.2

*Grain_1713:
XU_1713 in out fe_tanh Vc=0.5031490178859607 Qo=1.7740585213116075e-13 K=2.62 tau=9.37440425957272e-08 off=-0.2

*Grain_1714:
XU_1714 in out fe_tanh Vc=0.04599540370751182 Qo=1.621756874957734e-14 K=2.62 tau=9.501046611865559e-08 off=-0.2

*Grain_1715:
XU_1715 in out fe_tanh Vc=0.6266624325651053 Qo=2.2095557955157573e-13 K=2.62 tau=9.207250506127177e-08 off=-0.2

*Grain_1716:
XU_1716 in out fe_tanh Vc=0.21897662035745125 Qo=7.720920154935135e-14 K=2.62 tau=9.117704701258847e-08 off=-0.2

*Grain_1717:
XU_1717 in out fe_tanh Vc=0.3430438865861052 Qo=1.2095421208192996e-13 K=2.62 tau=1.1183410060823632e-07 off=-0.2

*Grain_1718:
XU_1718 in out fe_tanh Vc=0.329770064000405 Qo=1.1627398073268044e-13 K=2.62 tau=9.207210611604623e-08 off=-0.2

*Grain_1719:
XU_1719 in out fe_tanh Vc=0.9221961914259613 Qo=3.251581447171075e-13 K=2.62 tau=1.0124250809692614e-07 off=-0.2

*Grain_1720:
XU_1720 in out fe_tanh Vc=1.1732635118023678 Qo=4.1368224062175014e-13 K=2.62 tau=1.026975242272264e-07 off=-0.2

*Grain_1721:
XU_1721 in out fe_tanh Vc=0.23645885447692314 Qo=8.33732812372189e-14 K=2.62 tau=9.342534952035802e-08 off=-0.2

*Grain_1722:
XU_1722 in out fe_tanh Vc=0.47692230868177155 Qo=1.6815854858972787e-13 K=2.62 tau=8.906132582582805e-08 off=-0.2

*Grain_1723:
XU_1723 in out fe_tanh Vc=0.6034534716977662 Qo=2.1277230713449178e-13 K=2.62 tau=1.0194794096126147e-07 off=-0.2

*Grain_1724:
XU_1724 in out fe_tanh Vc=0.724872888006065 Qo=2.555837094223207e-13 K=2.62 tau=1.1411720070812349e-07 off=-0.2

*Grain_1725:
XU_1725 in out fe_tanh Vc=0.14549765363147876 Qo=5.1301173823273407e-14 K=2.62 tau=1.0093466805439865e-07 off=-0.2

*Grain_1726:
XU_1726 in out fe_tanh Vc=0.20260375048680587 Qo=7.143627379240442e-14 K=2.62 tau=8.83099309032778e-08 off=-0.2

*Grain_1727:
XU_1727 in out fe_tanh Vc=0.3493377743374918 Qo=1.2317338071798143e-13 K=2.62 tau=8.58019130568902e-08 off=-0.2

*Grain_1728:
XU_1728 in out fe_tanh Vc=0.381731965072927 Qo=1.3459528319066354e-13 K=2.62 tau=9.459752294012335e-08 off=-0.2

*Grain_1729:
XU_1729 in out fe_tanh Vc=0.22312932402312766 Qo=7.867340779097914e-14 K=2.62 tau=1.0417867320501366e-07 off=-0.2

*Grain_1730:
XU_1730 in out fe_tanh Vc=0.768779359169111 Qo=2.710647392044714e-13 K=2.62 tau=1.0548849198503456e-07 off=-0.2

*Grain_1731:
XU_1731 in out fe_tanh Vc=0.6462814280413886 Qo=2.2787306221913863e-13 K=2.62 tau=1.0858755094651522e-07 off=-0.2

*Grain_1732:
XU_1732 in out fe_tanh Vc=0.7467372615152688 Qo=2.632928923399617e-13 K=2.62 tau=1.0954713202489644e-07 off=-0.2

*Grain_1733:
XU_1733 in out fe_tanh Vc=0.525087214735055 Qo=1.8514106449943147e-13 K=2.62 tau=1.1253883530426605e-07 off=-0.2

*Grain_1734:
XU_1734 in out fe_tanh Vc=0.30843513846001896 Qo=1.0875147644250032e-13 K=2.62 tau=9.077104240623142e-08 off=-0.2

*Grain_1735:
XU_1735 in out fe_tanh Vc=0.5267871690275713 Qo=1.8574045320760185e-13 K=2.62 tau=8.695917943718849e-08 off=-0.2

*Grain_1736:
XU_1736 in out fe_tanh Vc=0.7109897017543907 Qo=2.5068862188419474e-13 K=2.62 tau=9.593354282003258e-08 off=-0.2

*Grain_1737:
XU_1737 in out fe_tanh Vc=0.6490835196178923 Qo=2.28861054694942e-13 K=2.62 tau=1.0554393520545267e-07 off=-0.2

*Grain_1738:
XU_1738 in out fe_tanh Vc=0.03881792013148139 Qo=1.3686852113553435e-14 K=2.62 tau=9.613491746674174e-08 off=-0.2

*Grain_1739:
XU_1739 in out fe_tanh Vc=0.2053911491773225 Qo=7.24190856877711e-14 K=2.62 tau=9.872407663202577e-08 off=-0.2

*Grain_1740:
XU_1740 in out fe_tanh Vc=0.2496708199903217 Qo=8.803170233496858e-14 K=2.62 tau=9.220846857235435e-08 off=-0.2

*Grain_1741:
XU_1741 in out fe_tanh Vc=0.49785094085496484 Qo=1.7553779746558776e-13 K=2.62 tau=1.1029136067316931e-07 off=-0.2

*Grain_1742:
XU_1742 in out fe_tanh Vc=0.6089502521808303 Qo=2.1471042286345253e-13 K=2.62 tau=1.0642648369683533e-07 off=-0.2

*Grain_1743:
XU_1743 in out fe_tanh Vc=0.5977473451535644 Qo=2.1076037785319127e-13 K=2.62 tau=1.115100368024817e-07 off=-0.2

*Grain_1744:
XU_1744 in out fe_tanh Vc=0.5757418749910774 Qo=2.0300144551516243e-13 K=2.62 tau=9.922444408435069e-08 off=-0.2

*Grain_1745:
XU_1745 in out fe_tanh Vc=0.20902488868286073 Qo=7.370030979929024e-14 K=2.62 tau=7.720283092476917e-08 off=-0.2

*Grain_1746:
XU_1746 in out fe_tanh Vc=0.73765839977674 Qo=2.6009176673730823e-13 K=2.62 tau=1.0574603418539566e-07 off=-0.2

*Grain_1747:
XU_1747 in out fe_tanh Vc=0.8502845497868172 Qo=2.998027418252459e-13 K=2.62 tau=9.707205984984172e-08 off=-0.2

*Grain_1748:
XU_1748 in out fe_tanh Vc=0.6063762773801911 Qo=2.1380286232643674e-13 K=2.62 tau=8.793155193420945e-08 off=-0.2

*Grain_1749:
XU_1749 in out fe_tanh Vc=-0.07460259676761799 Qo=2.6304209648196838e-14 K=2.62 tau=9.102985187768703e-08 off=-0.2

*Grain_1750:
XU_1750 in out fe_tanh Vc=0.7816246067667252 Qo=2.7559385883878016e-13 K=2.62 tau=8.605419003291942e-08 off=-0.2

*Grain_1751:
XU_1751 in out fe_tanh Vc=-0.2759819637207899 Qo=9.730877673662648e-14 K=2.62 tau=9.593630310586445e-08 off=-0.2

*Grain_1752:
XU_1752 in out fe_tanh Vc=0.4589800145850135 Qo=1.6183225586079182e-13 K=2.62 tau=9.089787325024933e-08 off=-0.2

*Grain_1753:
XU_1753 in out fe_tanh Vc=0.34184122956866 Qo=1.2053016595361228e-13 K=2.62 tau=9.616061463601814e-08 off=-0.2

*Grain_1754:
XU_1754 in out fe_tanh Vc=0.5323215432933299 Qo=1.8769182416874364e-13 K=2.62 tau=1.0675764815613124e-07 off=-0.2

*Grain_1755:
XU_1755 in out fe_tanh Vc=0.3526861302128176 Qo=1.24353981109087e-13 K=2.62 tau=9.273966275375104e-08 off=-0.2

*Grain_1756:
XU_1756 in out fe_tanh Vc=0.6542023526377752 Qo=2.306659095222951e-13 K=2.62 tau=1.2069665371262449e-07 off=-0.2

*Grain_1757:
XU_1757 in out fe_tanh Vc=0.15911674016641458 Qo=5.6103142158876755e-14 K=2.62 tau=1.1348431809853446e-07 off=-0.2

*Grain_1758:
XU_1758 in out fe_tanh Vc=0.5077689007343699 Qo=1.7903478158214485e-13 K=2.62 tau=1.0739017481181143e-07 off=-0.2

*Grain_1759:
XU_1759 in out fe_tanh Vc=0.1520802141410894 Qo=5.362212589691351e-14 K=2.62 tau=1.2141755004915196e-07 off=-0.2

*Grain_1760:
XU_1760 in out fe_tanh Vc=0.5749465468542997 Qo=2.027210199139722e-13 K=2.62 tau=9.640116030579413e-08 off=-0.2

*Grain_1761:
XU_1761 in out fe_tanh Vc=0.05197999198880793 Qo=1.8327681153569216e-14 K=2.62 tau=9.826193382392963e-08 off=-0.2

*Grain_1762:
XU_1762 in out fe_tanh Vc=0.2822728655026038 Qo=9.952689254646212e-14 K=2.62 tau=8.678449478837402e-08 off=-0.2

*Grain_1763:
XU_1763 in out fe_tanh Vc=0.12612605496265017 Qo=4.447092106152537e-14 K=2.62 tau=1.0722675730998602e-07 off=-0.2

*Grain_1764:
XU_1764 in out fe_tanh Vc=0.158735919368525 Qo=5.596886814510101e-14 K=2.62 tau=8.270908221378046e-08 off=-0.2

*Grain_1765:
XU_1765 in out fe_tanh Vc=0.44522984506928187 Qo=1.5698406883632832e-13 K=2.62 tau=1.0344748642205699e-07 off=-0.2

*Grain_1766:
XU_1766 in out fe_tanh Vc=0.8102480788052842 Qo=2.856862395598809e-13 K=2.62 tau=9.937387926984809e-08 off=-0.2

*Grain_1767:
XU_1767 in out fe_tanh Vc=0.09060299575663766 Qo=3.194580749730356e-14 K=2.62 tau=9.675717383574172e-08 off=-0.2

*Grain_1768:
XU_1768 in out fe_tanh Vc=0.5092021980971236 Qo=1.7954014943730844e-13 K=2.62 tau=8.766811837878043e-08 off=-0.2

*Grain_1769:
XU_1769 in out fe_tanh Vc=0.7166389030427669 Qo=2.5268047982845883e-13 K=2.62 tau=8.85104538263919e-08 off=-0.2

*Grain_1770:
XU_1770 in out fe_tanh Vc=0.18333877254207542 Qo=6.464361454617778e-14 K=2.62 tau=9.108388300582756e-08 off=-0.2

*Grain_1771:
XU_1771 in out fe_tanh Vc=0.34048685052367156 Qo=1.200526239927946e-13 K=2.62 tau=1.0135896864674817e-07 off=-0.2

*Grain_1772:
XU_1772 in out fe_tanh Vc=0.5564248050887005 Qo=1.9619041910969082e-13 K=2.62 tau=9.535399429970976e-08 off=-0.2

*Grain_1773:
XU_1773 in out fe_tanh Vc=-0.22358982088035056 Qo=7.883577487201332e-14 K=2.62 tau=9.490339883332254e-08 off=-0.2

*Grain_1774:
XU_1774 in out fe_tanh Vc=0.6074608345410875 Qo=2.141852674996043e-13 K=2.62 tau=1.0643360407733096e-07 off=-0.2

*Grain_1775:
XU_1775 in out fe_tanh Vc=0.4235634785930285 Qo=1.49344701430911e-13 K=2.62 tau=9.697266232016633e-08 off=-0.2

*Grain_1776:
XU_1776 in out fe_tanh Vc=0.580006157299795 Qo=2.0450499339027192e-13 K=2.62 tau=9.42156155203136e-08 off=-0.2

*Grain_1777:
XU_1777 in out fe_tanh Vc=0.153466800214986 Qo=5.411102376861437e-14 K=2.62 tau=9.823794686900865e-08 off=-0.2

*Grain_1778:
XU_1778 in out fe_tanh Vc=-0.004950909531755865 Qo=1.745646504480523e-15 K=2.62 tau=1.0453331979842795e-07 off=-0.2

*Grain_1779:
XU_1779 in out fe_tanh Vc=0.3315996267137123 Qo=1.1691906821301661e-13 K=2.62 tau=9.875982320683018e-08 off=-0.2

*Grain_1780:
XU_1780 in out fe_tanh Vc=0.5973790623620601 Qo=2.1063052462854108e-13 K=2.62 tau=9.937969624427609e-08 off=-0.2

*Grain_1781:
XU_1781 in out fe_tanh Vc=0.22310278374044895 Qo=7.866404992422984e-14 K=2.62 tau=9.828841279961317e-08 off=-0.2

*Grain_1782:
XU_1782 in out fe_tanh Vc=0.5713613525659975 Qo=2.0145691241269079e-13 K=2.62 tau=1.0065004758509016e-07 off=-0.2

*Grain_1783:
XU_1783 in out fe_tanh Vc=0.34655875023963706 Qo=1.2219352162922794e-13 K=2.62 tau=8.865261149684054e-08 off=-0.2

*Grain_1784:
XU_1784 in out fe_tanh Vc=-0.17485663906925059 Qo=6.165289000306082e-14 K=2.62 tau=8.411867994860248e-08 off=-0.2

*Grain_1785:
XU_1785 in out fe_tanh Vc=0.30827799795062205 Qo=1.086960701016691e-13 K=2.62 tau=1.0645761274781668e-07 off=-0.2

*Grain_1786:
XU_1786 in out fe_tanh Vc=-0.12689523286283627 Qo=4.474212632273468e-14 K=2.62 tau=9.877948545933898e-08 off=-0.2

*Grain_1787:
XU_1787 in out fe_tanh Vc=0.3888921611075543 Qo=1.3711990439391338e-13 K=2.62 tau=9.181775732679841e-08 off=-0.2

*Grain_1788:
XU_1788 in out fe_tanh Vc=0.5244056136140068 Qo=1.849007380287545e-13 K=2.62 tau=1.0316765608499302e-07 off=-0.2

*Grain_1789:
XU_1789 in out fe_tanh Vc=0.8750604322051004 Qo=3.0853849679339574e-13 K=2.62 tau=1.0307063681434424e-07 off=-0.2

*Grain_1790:
XU_1790 in out fe_tanh Vc=0.4706434803580888 Qo=1.6594468977345036e-13 K=2.62 tau=9.827304283453002e-08 off=-0.2

*Grain_1791:
XU_1791 in out fe_tanh Vc=0.5437880460255948 Qo=1.9173481067148745e-13 K=2.62 tau=1.0750365728605457e-07 off=-0.2

*Grain_1792:
XU_1792 in out fe_tanh Vc=0.7013199446523117 Qo=2.472791518512343e-13 K=2.62 tau=1.0437104693568986e-07 off=-0.2

*Grain_1793:
XU_1793 in out fe_tanh Vc=0.883281052343878 Qo=3.114370140694385e-13 K=2.62 tau=9.415830843079433e-08 off=-0.2

*Grain_1794:
XU_1794 in out fe_tanh Vc=0.4282475336809534 Qo=1.5099625744068734e-13 K=2.62 tau=1.0364498753891492e-07 off=-0.2

*Grain_1795:
XU_1795 in out fe_tanh Vc=-0.07858170377304713 Qo=2.770720725710646e-14 K=2.62 tau=8.868051788530389e-08 off=-0.2

*Grain_1796:
XU_1796 in out fe_tanh Vc=0.2791053665214245 Qo=9.8410060681736e-14 K=2.62 tau=1.018107556227504e-07 off=-0.2

*Grain_1797:
XU_1797 in out fe_tanh Vc=0.7682177952433782 Qo=2.7086673677729913e-13 K=2.62 tau=1.0613432592259909e-07 off=-0.2

*Grain_1798:
XU_1798 in out fe_tanh Vc=0.40967822079044147 Qo=1.4444888348242576e-13 K=2.62 tau=9.140818741160785e-08 off=-0.2

*Grain_1799:
XU_1799 in out fe_tanh Vc=0.1889286345633846 Qo=6.661454999459146e-14 K=2.62 tau=1.1911389331344835e-07 off=-0.2

*Grain_1800:
XU_1800 in out fe_tanh Vc=0.059289532994819316 Qo=2.0904960060537137e-14 K=2.62 tau=8.971074776689602e-08 off=-0.2

*Grain_1801:
XU_1801 in out fe_tanh Vc=0.28651015122441503 Qo=1.0102092166602508e-13 K=2.62 tau=1.0566053649439984e-07 off=-0.2

*Grain_1802:
XU_1802 in out fe_tanh Vc=0.6325361242722798 Qo=2.2302659081349813e-13 K=2.62 tau=1.1072275659050573e-07 off=-0.2

*Grain_1803:
XU_1803 in out fe_tanh Vc=0.7903825715511668 Qo=2.786818390400467e-13 K=2.62 tau=8.580250194021113e-08 off=-0.2

*Grain_1804:
XU_1804 in out fe_tanh Vc=0.9311321820606555 Qo=3.2830889524394903e-13 K=2.62 tau=1.2399224185659692e-07 off=-0.2

*Grain_1805:
XU_1805 in out fe_tanh Vc=0.5664857861806483 Qo=1.9973783122905033e-13 K=2.62 tau=1.1012635606330733e-07 off=-0.2

*Grain_1806:
XU_1806 in out fe_tanh Vc=0.6760957721850409 Qo=2.383853338136648e-13 K=2.62 tau=9.787757643304707e-08 off=-0.2

*Grain_1807:
XU_1807 in out fe_tanh Vc=0.34269723479861725 Qo=1.208319857561975e-13 K=2.62 tau=1.0398572985262936e-07 off=-0.2

*Grain_1808:
XU_1808 in out fe_tanh Vc=0.05161725920043897 Qo=1.8199784810480076e-14 K=2.62 tau=8.95055891566477e-08 off=-0.2

*Grain_1809:
XU_1809 in out fe_tanh Vc=-0.6687634970710883 Qo=2.358000390631825e-13 K=2.62 tau=1.1000087443607249e-07 off=-0.2

*Grain_1810:
XU_1810 in out fe_tanh Vc=0.35740323751013564 Qo=1.2601719103284063e-13 K=2.62 tau=1.0632641177123778e-07 off=-0.2

*Grain_1811:
XU_1811 in out fe_tanh Vc=0.38252187087438516 Qo=1.348737969248249e-13 K=2.62 tau=9.752423621094174e-08 off=-0.2

*Grain_1812:
XU_1812 in out fe_tanh Vc=0.3931439158150291 Qo=1.3861903514865767e-13 K=2.62 tau=8.417669990630566e-08 off=-0.2

*Grain_1813:
XU_1813 in out fe_tanh Vc=0.2479615417689622 Qo=8.74290260927221e-14 K=2.62 tau=8.690664329182825e-08 off=-0.2

*Grain_1814:
XU_1814 in out fe_tanh Vc=0.126370706949904 Qo=4.455718316824021e-14 K=2.62 tau=8.650112086912195e-08 off=-0.2

*Grain_1815:
XU_1815 in out fe_tanh Vc=0.10929420016756919 Qo=3.8536159317548154e-14 K=2.62 tau=9.825910564131092e-08 off=-0.2

*Grain_1816:
XU_1816 in out fe_tanh Vc=0.5131322012147718 Qo=1.8092583345373338e-13 K=2.62 tau=1.0509365373286416e-07 off=-0.2

*Grain_1817:
XU_1817 in out fe_tanh Vc=-0.04720410079359327 Qo=1.66437445521769e-14 K=2.62 tau=1.0594758450902542e-07 off=-0.2

*Grain_1818:
XU_1818 in out fe_tanh Vc=0.545742274367897 Qo=1.9242385413972605e-13 K=2.62 tau=1.1035966816227545e-07 off=-0.2

*Grain_1819:
XU_1819 in out fe_tanh Vc=0.8506558879706487 Qo=2.999336723539554e-13 K=2.62 tau=1.060988003843871e-07 off=-0.2

*Grain_1820:
XU_1820 in out fe_tanh Vc=0.5260236517498059 Qo=1.854712438313261e-13 K=2.62 tau=8.72720719105261e-08 off=-0.2

*Grain_1821:
XU_1821 in out fe_tanh Vc=0.4910121491597878 Qo=1.7312650056327447e-13 K=2.62 tau=9.595704349283934e-08 off=-0.2

*Grain_1822:
XU_1822 in out fe_tanh Vc=0.45076442281985485 Qo=1.5893551154439915e-13 K=2.62 tau=8.534335484370618e-08 off=-0.2

*Grain_1823:
XU_1823 in out fe_tanh Vc=0.2257824452732173 Qo=7.960887465953643e-14 K=2.62 tau=1.0744655622126019e-07 off=-0.2

*Grain_1824:
XU_1824 in out fe_tanh Vc=1.010973579515277 Qo=3.564602592479829e-13 K=2.62 tau=1.0301975718386658e-07 off=-0.2

*Grain_1825:
XU_1825 in out fe_tanh Vc=0.7057369241256282 Qo=2.4883653938346466e-13 K=2.62 tau=1.2165788658799264e-07 off=-0.2

*Grain_1826:
XU_1826 in out fe_tanh Vc=0.5832783051987774 Qo=2.05658723529222e-13 K=2.62 tau=1.0630937336521192e-07 off=-0.2

*Grain_1827:
XU_1827 in out fe_tanh Vc=0.7567973658510312 Qo=2.6683999532291695e-13 K=2.62 tau=1.0047945300298117e-07 off=-0.2

*Grain_1828:
XU_1828 in out fe_tanh Vc=0.48796127110026344 Qo=1.720507881944572e-13 K=2.62 tau=1.1577827373658904e-07 off=-0.2

*Grain_1829:
XU_1829 in out fe_tanh Vc=0.4962659573454017 Qo=1.7497894642915063e-13 K=2.62 tau=9.087301205045307e-08 off=-0.2

*Grain_1830:
XU_1830 in out fe_tanh Vc=-0.043880913289727264 Qo=1.547201830417179e-14 K=2.62 tau=7.899109054277776e-08 off=-0.2

*Grain_1831:
XU_1831 in out fe_tanh Vc=0.9112413504312364 Qo=3.212955655754525e-13 K=2.62 tau=1.0612698449189157e-07 off=-0.2

*Grain_1832:
XU_1832 in out fe_tanh Vc=0.47275750892025425 Qo=1.6669007737268755e-13 K=2.62 tau=1.0245161546105716e-07 off=-0.2

*Grain_1833:
XU_1833 in out fe_tanh Vc=0.3745413781751208 Qo=1.320599464403539e-13 K=2.62 tau=1.0540425135891275e-07 off=-0.2

*Grain_1834:
XU_1834 in out fe_tanh Vc=0.25462033441591536 Qo=8.977685693747032e-14 K=2.62 tau=1.062669724084104e-07 off=-0.2

*Grain_1835:
XU_1835 in out fe_tanh Vc=0.021252998377423282 Qo=7.493617503877393e-15 K=2.62 tau=9.77210408647206e-08 off=-0.2

*Grain_1836:
XU_1836 in out fe_tanh Vc=0.3842265543951208 Qo=1.3547485311664797e-13 K=2.62 tau=1.0368031286104999e-07 off=-0.2

*Grain_1837:
XU_1837 in out fe_tanh Vc=1.1169249130120065 Qo=3.9381775361892553e-13 K=2.62 tau=1.1007141035960179e-07 off=-0.2

*Grain_1838:
XU_1838 in out fe_tanh Vc=0.1236717305465529 Qo=4.3605548181988636e-14 K=2.62 tau=1.1521652379245177e-07 off=-0.2

*Grain_1839:
XU_1839 in out fe_tanh Vc=0.9408262505008325 Qo=3.3172693723769725e-13 K=2.62 tau=9.411964430932549e-08 off=-0.2

*Grain_1840:
XU_1840 in out fe_tanh Vc=0.509946966777232 Qo=1.7980274822541768e-13 K=2.62 tau=9.306568069694727e-08 off=-0.2

*Grain_1841:
XU_1841 in out fe_tanh Vc=0.20647154221335048 Qo=7.280002262768293e-14 K=2.62 tau=1.0729567904930217e-07 off=-0.2

*Grain_1842:
XU_1842 in out fe_tanh Vc=0.5152074789016676 Qo=1.8165755784027682e-13 K=2.62 tau=1.0514477384226483e-07 off=-0.2

*Grain_1843:
XU_1843 in out fe_tanh Vc=0.30355466348163307 Qo=1.070306645327738e-13 K=2.62 tau=1.0106644459861055e-07 off=-0.2

*Grain_1844:
XU_1844 in out fe_tanh Vc=0.657621469120389 Qo=2.318714594718555e-13 K=2.62 tau=1.1165092542580459e-07 off=-0.2

*Grain_1845:
XU_1845 in out fe_tanh Vc=-0.05687101624976626 Qo=2.005221264615807e-14 K=2.62 tau=1.082259707306653e-07 off=-0.2

*Grain_1846:
XU_1846 in out fe_tanh Vc=0.4900226041248997 Qo=1.7277759581757093e-13 K=2.62 tau=1.1067526087991162e-07 off=-0.2

*Grain_1847:
XU_1847 in out fe_tanh Vc=0.5658079157903039 Qo=1.9949882018071556e-13 K=2.62 tau=1.0563006623168978e-07 off=-0.2

*Grain_1848:
XU_1848 in out fe_tanh Vc=0.6261789348665112 Qo=2.2078510257920096e-13 K=2.62 tau=9.609559116230835e-08 off=-0.2

*Grain_1849:
XU_1849 in out fe_tanh Vc=0.1638864615930679 Qo=5.778490335495142e-14 K=2.62 tau=8.971502576265157e-08 off=-0.2

*Grain_1850:
XU_1850 in out fe_tanh Vc=-0.011915252717785207 Qo=4.201211741679117e-15 K=2.62 tau=1.1297280877129642e-07 off=-0.2

*Grain_1851:
XU_1851 in out fe_tanh Vc=0.8577648757290646 Qo=3.024402379761457e-13 K=2.62 tau=1.0078883126819881e-07 off=-0.2

*Grain_1852:
XU_1852 in out fe_tanh Vc=-0.0037974003894867825 Qo=1.33892947821036e-15 K=2.62 tau=1.0667011815025346e-07 off=-0.2

*Grain_1853:
XU_1853 in out fe_tanh Vc=0.35568464137049377 Qo=1.2541122937578818e-13 K=2.62 tau=9.601193824589773e-08 off=-0.2

*Grain_1854:
XU_1854 in out fe_tanh Vc=0.6434754649508196 Qo=2.2688370468203657e-13 K=2.62 tau=1.1542987097482744e-07 off=-0.2

*Grain_1855:
XU_1855 in out fe_tanh Vc=0.5734251086448119 Qo=2.021845743830773e-13 K=2.62 tau=8.637670370647623e-08 off=-0.2

*Grain_1856:
XU_1856 in out fe_tanh Vc=0.9334406666357773 Qo=3.291228462974597e-13 K=2.62 tau=9.97533847156899e-08 off=-0.2

*Grain_1857:
XU_1857 in out fe_tanh Vc=0.7673591391174294 Qo=2.705639822924517e-13 K=2.62 tau=9.706274449618492e-08 off=-0.2

*Grain_1858:
XU_1858 in out fe_tanh Vc=0.677546448016783 Qo=2.388968291618572e-13 K=2.62 tau=9.274373769142119e-08 off=-0.2

*Grain_1859:
XU_1859 in out fe_tanh Vc=-0.13700008800311964 Qo=4.830500803987681e-14 K=2.62 tau=1.0417972998435477e-07 off=-0.2

*Grain_1860:
XU_1860 in out fe_tanh Vc=1.036004423164755 Qo=3.652859112702312e-13 K=2.62 tau=9.857997317096194e-08 off=-0.2

*Grain_1861:
XU_1861 in out fe_tanh Vc=0.3424145731746206 Qo=1.207323217908765e-13 K=2.62 tau=1.0334616078199157e-07 off=-0.2

*Grain_1862:
XU_1862 in out fe_tanh Vc=0.13662234728791323 Qo=4.8171820035759486e-14 K=2.62 tau=9.980213045013328e-08 off=-0.2

*Grain_1863:
XU_1863 in out fe_tanh Vc=0.5581803555247088 Qo=1.968094105217537e-13 K=2.62 tau=1.0564465868380105e-07 off=-0.2

*Grain_1864:
XU_1864 in out fe_tanh Vc=0.3248326795266092 Qo=1.145331030428994e-13 K=2.62 tau=1.0726495459961024e-07 off=-0.2

*Grain_1865:
XU_1865 in out fe_tanh Vc=0.5632871020979584 Qo=1.9861000377591877e-13 K=2.62 tau=9.726138485925249e-08 off=-0.2

*Grain_1866:
XU_1866 in out fe_tanh Vc=-0.023933310664424057 Qo=8.438671689317076e-15 K=2.62 tau=1.139190225382132e-07 off=-0.2

*Grain_1867:
XU_1867 in out fe_tanh Vc=0.21262696797142125 Qo=7.497037080093155e-14 K=2.62 tau=8.776353419848425e-08 off=-0.2

*Grain_1868:
XU_1868 in out fe_tanh Vc=0.4231162971613631 Qo=1.4918702925006254e-13 K=2.62 tau=9.531882543712691e-08 off=-0.2

*Grain_1869:
XU_1869 in out fe_tanh Vc=0.09032187957775278 Qo=3.1846688442132854e-14 K=2.62 tau=1.0149306557996131e-07 off=-0.2

*Grain_1870:
XU_1870 in out fe_tanh Vc=0.13158547497364192 Qo=4.639586382154765e-14 K=2.62 tau=1.0071930003487112e-07 off=-0.2

*Grain_1871:
XU_1871 in out fe_tanh Vc=0.12595673436350757 Qo=4.4411220129780605e-14 K=2.62 tau=1.0305272097040441e-07 off=-0.2

*Grain_1872:
XU_1872 in out fe_tanh Vc=0.22063717380022085 Qo=7.779469786962966e-14 K=2.62 tau=1.1932512564764763e-07 off=-0.2

*Grain_1873:
XU_1873 in out fe_tanh Vc=0.278568703212077 Qo=9.822083798961519e-14 K=2.62 tau=9.687627672745615e-08 off=-0.2

*Grain_1874:
XU_1874 in out fe_tanh Vc=0.5516497571461279 Qo=1.9450677983165243e-13 K=2.62 tau=1.0374439803226299e-07 off=-0.2

*Grain_1875:
XU_1875 in out fe_tanh Vc=0.6730245798905001 Qo=2.3730245882692445e-13 K=2.62 tau=9.120748353428285e-08 off=-0.2

*Grain_1876:
XU_1876 in out fe_tanh Vc=0.7361654495231833 Qo=2.595653658053647e-13 K=2.62 tau=1.0550145395701734e-07 off=-0.2

*Grain_1877:
XU_1877 in out fe_tanh Vc=0.00017891825926696914 Qo=6.308498102698231e-17 K=2.62 tau=1.2110309421736617e-07 off=-0.2

*Grain_1878:
XU_1878 in out fe_tanh Vc=0.8644399473865876 Qo=3.047938086546993e-13 K=2.62 tau=1.0152150598725313e-07 off=-0.2

*Grain_1879:
XU_1879 in out fe_tanh Vc=0.6815813455736659 Qo=2.403194980211712e-13 K=2.62 tau=1.1127173083193182e-07 off=-0.2

*Grain_1880:
XU_1880 in out fe_tanh Vc=1.0542018587196689 Qo=3.717021645996834e-13 K=2.62 tau=9.723963159956801e-08 off=-0.2

*Grain_1881:
XU_1881 in out fe_tanh Vc=0.43184171670469845 Qo=1.5226353428984411e-13 K=2.62 tau=7.908867362579091e-08 off=-0.2

*Grain_1882:
XU_1882 in out fe_tanh Vc=0.24003029252691704 Qo=8.463253841167379e-14 K=2.62 tau=9.528507688073235e-08 off=-0.2

*Grain_1883:
XU_1883 in out fe_tanh Vc=0.6328011080837239 Qo=2.2312002173992172e-13 K=2.62 tau=9.224128763473454e-08 off=-0.2

*Grain_1884:
XU_1884 in out fe_tanh Vc=0.5908569355389032 Qo=2.0833088093325734e-13 K=2.62 tau=1.0258861694404636e-07 off=-0.2

*Grain_1885:
XU_1885 in out fe_tanh Vc=-0.07480745783962456 Qo=2.637644183340616e-14 K=2.62 tau=1.1541403074265118e-07 off=-0.2

*Grain_1886:
XU_1886 in out fe_tanh Vc=0.752048307239932 Qo=2.651655196511512e-13 K=2.62 tau=1.0762287400263769e-07 off=-0.2

*Grain_1887:
XU_1887 in out fe_tanh Vc=0.4007583552877587 Qo=1.4130381853318356e-13 K=2.62 tau=9.386621815528529e-08 off=-0.2

*Grain_1888:
XU_1888 in out fe_tanh Vc=0.26524192036994365 Qo=9.352193332671976e-14 K=2.62 tau=1.0957858005428014e-07 off=-0.2

*Grain_1889:
XU_1889 in out fe_tanh Vc=0.23272850118442037 Qo=8.205799196688047e-14 K=2.62 tau=1.0155257805373225e-07 off=-0.2

*Grain_1890:
XU_1890 in out fe_tanh Vc=0.19497740671952396 Qo=6.874729305988819e-14 K=2.62 tau=1.0601817594599775e-07 off=-0.2

*Grain_1891:
XU_1891 in out fe_tanh Vc=0.5324540522480248 Qo=1.8773854564327105e-13 K=2.62 tau=7.261920082060084e-08 off=-0.2

*Grain_1892:
XU_1892 in out fe_tanh Vc=0.11250377782012988 Qo=3.966782774617006e-14 K=2.62 tau=9.832595619705691e-08 off=-0.2

*Grain_1893:
XU_1893 in out fe_tanh Vc=0.8061950983004382 Qo=2.8425719481454034e-13 K=2.62 tau=1.0806332146698859e-07 off=-0.2

*Grain_1894:
XU_1894 in out fe_tanh Vc=0.5733593709427497 Qo=2.0216139585616594e-13 K=2.62 tau=1.0134616268886151e-07 off=-0.2

*Grain_1895:
XU_1895 in out fe_tanh Vc=0.5753394111627285 Qo=2.0285954036205248e-13 K=2.62 tau=1.0776307707042168e-07 off=-0.2

*Grain_1896:
XU_1896 in out fe_tanh Vc=0.018095692370433625 Qo=6.3803795908585795e-15 K=2.62 tau=9.734592393729195e-08 off=-0.2

*Grain_1897:
XU_1897 in out fe_tanh Vc=0.3104102627787575 Qo=1.0944788764549346e-13 K=2.62 tau=1.1094787098356195e-07 off=-0.2

*Grain_1898:
XU_1898 in out fe_tanh Vc=0.3815653662643215 Qo=1.3453654193796494e-13 K=2.62 tau=1.0802884604871132e-07 off=-0.2

*Grain_1899:
XU_1899 in out fe_tanh Vc=0.21036467934791978 Qo=7.417270802757427e-14 K=2.62 tau=9.139979664232573e-08 off=-0.2

*Grain_1900:
XU_1900 in out fe_tanh Vc=0.14652385014330083 Qo=5.166300155255873e-14 K=2.62 tau=1.1012299443239112e-07 off=-0.2

*Grain_1901:
XU_1901 in out fe_tanh Vc=0.5136880943095978 Qo=1.81121836396551e-13 K=2.62 tau=9.780055255431422e-08 off=-0.2

*Grain_1902:
XU_1902 in out fe_tanh Vc=0.4311636140119239 Qo=1.520244413337462e-13 K=2.62 tau=1.076743956400441e-07 off=-0.2

*Grain_1903:
XU_1903 in out fe_tanh Vc=0.7323016643662581 Qo=2.582030296507676e-13 K=2.62 tau=7.526260648326915e-08 off=-0.2

*Grain_1904:
XU_1904 in out fe_tanh Vc=0.2060118889794968 Qo=7.263795300071778e-14 K=2.62 tau=9.325105604773378e-08 off=-0.2

*Grain_1905:
XU_1905 in out fe_tanh Vc=0.6833640648308796 Qo=2.40948068917057e-13 K=2.62 tau=9.905265413624036e-08 off=-0.2

*Grain_1906:
XU_1906 in out fe_tanh Vc=-0.25163574948021733 Qo=8.872451893232023e-14 K=2.62 tau=1.122709388663158e-07 off=-0.2

*Grain_1907:
XU_1907 in out fe_tanh Vc=-0.3553101273616594 Qo=1.2527917907953306e-13 K=2.62 tau=1.1597408548529099e-07 off=-0.2

*Grain_1908:
XU_1908 in out fe_tanh Vc=0.7107325787868641 Qo=2.505979626211633e-13 K=2.62 tau=9.613606683951643e-08 off=-0.2

*Grain_1909:
XU_1909 in out fe_tanh Vc=0.24127633192747883 Qo=8.507188078100693e-14 K=2.62 tau=1.1425175977518482e-07 off=-0.2

*Grain_1910:
XU_1910 in out fe_tanh Vc=0.3832255916532946 Qo=1.3512192258940312e-13 K=2.62 tau=9.222168628059374e-08 off=-0.2

*Grain_1911:
XU_1911 in out fe_tanh Vc=0.20906472654102326 Qo=7.371435627244863e-14 K=2.62 tau=1.092454578829199e-07 off=-0.2

*Grain_1912:
XU_1912 in out fe_tanh Vc=0.4245595294507012 Qo=1.4969590007165135e-13 K=2.62 tau=1.0794207482750197e-07 off=-0.2

*Grain_1913:
XU_1913 in out fe_tanh Vc=0.0001670930786541458 Qo=5.891552790544549e-17 K=2.62 tau=8.857276453866948e-08 off=-0.2

*Grain_1914:
XU_1914 in out fe_tanh Vc=0.7968147082083168 Qo=2.809497530061322e-13 K=2.62 tau=1.100369966745292e-07 off=-0.2

*Grain_1915:
XU_1915 in out fe_tanh Vc=0.5720492371506647 Qo=2.0169945437654777e-13 K=2.62 tau=1.1486802916984495e-07 off=-0.2

*Grain_1916:
XU_1916 in out fe_tanh Vc=0.9252505288762678 Qo=3.2623507683623283e-13 K=2.62 tau=9.974804346014425e-08 off=-0.2

*Grain_1917:
XU_1917 in out fe_tanh Vc=0.8285408270463341 Qo=2.9213609929161505e-13 K=2.62 tau=1.0750043958421331e-07 off=-0.2

*Grain_1918:
XU_1918 in out fe_tanh Vc=0.5161116263018862 Qo=1.8197635214233449e-13 K=2.62 tau=8.433518283791737e-08 off=-0.2

*Grain_1919:
XU_1919 in out fe_tanh Vc=0.17510729208429898 Qo=6.174126801860529e-14 K=2.62 tau=9.924925183747655e-08 off=-0.2

*Grain_1920:
XU_1920 in out fe_tanh Vc=0.8408839389729688 Qo=2.964881703708658e-13 K=2.62 tau=1.0646259958099786e-07 off=-0.2

*Grain_1921:
XU_1921 in out fe_tanh Vc=0.16926075028766557 Qo=5.967982957277435e-14 K=2.62 tau=1.0221489805232365e-07 off=-0.2

*Grain_1922:
XU_1922 in out fe_tanh Vc=0.9163013792442156 Qo=3.230796865643923e-13 K=2.62 tau=1.1361219334961209e-07 off=-0.2

*Grain_1923:
XU_1923 in out fe_tanh Vc=0.31970751126112773 Qo=1.1272601446450252e-13 K=2.62 tau=9.696256130972749e-08 off=-0.2

*Grain_1924:
XU_1924 in out fe_tanh Vc=0.03815538095228088 Qo=1.3453246713407377e-14 K=2.62 tau=9.746932596440428e-08 off=-0.2

*Grain_1925:
XU_1925 in out fe_tanh Vc=0.30429688052438836 Qo=1.0729236363633066e-13 K=2.62 tau=9.002200215729766e-08 off=-0.2

*Grain_1926:
XU_1926 in out fe_tanh Vc=0.8001184372094553 Qo=2.821146183597803e-13 K=2.62 tau=1.0146048913794263e-07 off=-0.2

*Grain_1927:
XU_1927 in out fe_tanh Vc=0.8948644395091967 Qo=3.1552121297985805e-13 K=2.62 tau=9.051288359209021e-08 off=-0.2

*Grain_1928:
XU_1928 in out fe_tanh Vc=-0.13174223586527162 Qo=4.645113631254297e-14 K=2.62 tau=1.1077374248882408e-07 off=-0.2

*Grain_1929:
XU_1929 in out fe_tanh Vc=0.569138343454464 Qo=2.00673099244608e-13 K=2.62 tau=9.333493515895841e-08 off=-0.2

*Grain_1930:
XU_1930 in out fe_tanh Vc=0.7606120663720424 Qo=2.681850246730658e-13 K=2.62 tau=8.662488856136682e-08 off=-0.2

*Grain_1931:
XU_1931 in out fe_tanh Vc=0.4188224306851455 Qo=1.476730502615883e-13 K=2.62 tau=9.28638207750222e-08 off=-0.2

*Grain_1932:
XU_1932 in out fe_tanh Vc=0.8212212501493124 Qo=2.895552818190665e-13 K=2.62 tau=7.49923449769242e-08 off=-0.2

*Grain_1933:
XU_1933 in out fe_tanh Vc=0.5706379608533034 Qo=2.0120185095246111e-13 K=2.62 tau=1.0095853656063231e-07 off=-0.2

*Grain_1934:
XU_1934 in out fe_tanh Vc=0.413311263634938 Qo=1.4572986195748066e-13 K=2.62 tau=1.1039228503613046e-07 off=-0.2

*Grain_1935:
XU_1935 in out fe_tanh Vc=-0.0839656533333652 Qo=2.960553980994054e-14 K=2.62 tau=1.1209427025705801e-07 off=-0.2

*Grain_1936:
XU_1936 in out fe_tanh Vc=0.33329017289296625 Qo=1.175151397044363e-13 K=2.62 tau=8.141566939733726e-08 off=-0.2

*Grain_1937:
XU_1937 in out fe_tanh Vc=0.4017360699664393 Qo=1.4164855200089705e-13 K=2.62 tau=1.0052054238565207e-07 off=-0.2

*Grain_1938:
XU_1938 in out fe_tanh Vc=-0.18374539254980454 Qo=6.478698513103524e-14 K=2.62 tau=1.0206775919282922e-07 off=-0.2

*Grain_1939:
XU_1939 in out fe_tanh Vc=0.2502496245732949 Qo=8.823578366397767e-14 K=2.62 tau=8.523777828838435e-08 off=-0.2

*Grain_1940:
XU_1940 in out fe_tanh Vc=0.6955966575041624 Qo=2.452611718941734e-13 K=2.62 tau=9.731043244775925e-08 off=-0.2

*Grain_1941:
XU_1941 in out fe_tanh Vc=0.26142028149481333 Qo=9.217445757484671e-14 K=2.62 tau=9.957545763553093e-08 off=-0.2

*Grain_1942:
XU_1942 in out fe_tanh Vc=0.7443405337321094 Qo=2.624478275190378e-13 K=2.62 tau=1.1642537284247301e-07 off=-0.2

*Grain_1943:
XU_1943 in out fe_tanh Vc=0.7732700835685291 Qo=2.7264812853932947e-13 K=2.62 tau=9.801932412607381e-08 off=-0.2

*Grain_1944:
XU_1944 in out fe_tanh Vc=0.38064370032025785 Qo=1.342115707537343e-13 K=2.62 tau=1.018473539305742e-07 off=-0.2

*Grain_1945:
XU_1945 in out fe_tanh Vc=0.4758201882271062 Qo=1.6776995075596364e-13 K=2.62 tau=9.162322007630314e-08 off=-0.2

*Grain_1946:
XU_1946 in out fe_tanh Vc=0.37247585590901106 Qo=1.3133166172809373e-13 K=2.62 tau=1.164968511285597e-07 off=-0.2

*Grain_1947:
XU_1947 in out fe_tanh Vc=0.6345280049697695 Qo=2.2372891016605593e-13 K=2.62 tau=1.022623195880342e-07 off=-0.2

*Grain_1948:
XU_1948 in out fe_tanh Vc=0.6324986058456639 Qo=2.2301336215119766e-13 K=2.62 tau=1.1502201974853797e-07 off=-0.2

*Grain_1949:
XU_1949 in out fe_tanh Vc=0.25773786427330736 Qo=9.087607013521985e-14 K=2.62 tau=1.0827300579912423e-07 off=-0.2

*Grain_1950:
XU_1950 in out fe_tanh Vc=0.5898693949370528 Qo=2.0798268293274949e-13 K=2.62 tau=8.455289303504147e-08 off=-0.2

*Grain_1951:
XU_1951 in out fe_tanh Vc=0.4985029057560964 Qo=1.7576767446968253e-13 K=2.62 tau=8.947973859382501e-08 off=-0.2

*Grain_1952:
XU_1952 in out fe_tanh Vc=0.425208964506767 Qo=1.499248850749597e-13 K=2.62 tau=9.82011059185956e-08 off=-0.2

*Grain_1953:
XU_1953 in out fe_tanh Vc=0.4383151801286032 Qo=1.5454601970496622e-13 K=2.62 tau=1.1031120624218864e-07 off=-0.2

*Grain_1954:
XU_1954 in out fe_tanh Vc=0.3838500439931687 Qo=1.3534209891000118e-13 K=2.62 tau=9.397275886014717e-08 off=-0.2

*Grain_1955:
XU_1955 in out fe_tanh Vc=0.45996203989116974 Qo=1.621785092172726e-13 K=2.62 tau=9.357294308314869e-08 off=-0.2

*Grain_1956:
XU_1956 in out fe_tanh Vc=0.409454903962443 Qo=1.4437014396240692e-13 K=2.62 tau=8.554661824867655e-08 off=-0.2

*Grain_1957:
XU_1957 in out fe_tanh Vc=0.37062321011329874 Qo=1.3067843535896255e-13 K=2.62 tau=1.0860972527629868e-07 off=-0.2

*Grain_1958:
XU_1958 in out fe_tanh Vc=0.27371384406620214 Qo=9.650905799376136e-14 K=2.62 tau=8.759016939753515e-08 off=-0.2

*Grain_1959:
XU_1959 in out fe_tanh Vc=0.6415680091203843 Qo=2.2621115278394732e-13 K=2.62 tau=9.300735237072117e-08 off=-0.2

*Grain_1960:
XU_1960 in out fe_tanh Vc=0.5886278819312967 Qo=2.07544936529818e-13 K=2.62 tau=9.79216454529547e-08 off=-0.2

*Grain_1961:
XU_1961 in out fe_tanh Vc=0.5526200192568261 Qo=1.9484888559042393e-13 K=2.62 tau=8.537851852474511e-08 off=-0.2

*Grain_1962:
XU_1962 in out fe_tanh Vc=0.41359911096815116 Qo=1.4583135435757898e-13 K=2.62 tau=1.1254024149147127e-07 off=-0.2

*Grain_1963:
XU_1963 in out fe_tanh Vc=0.8490823792682451 Qo=2.993788672320879e-13 K=2.62 tau=1.0097871831187301e-07 off=-0.2

*Grain_1964:
XU_1964 in out fe_tanh Vc=0.23005702998034247 Qo=8.111605506835566e-14 K=2.62 tau=1.1765638233433558e-07 off=-0.2

*Grain_1965:
XU_1965 in out fe_tanh Vc=0.6697784734312594 Qo=2.361579106671572e-13 K=2.62 tau=1.0520663954158783e-07 off=-0.2

*Grain_1966:
XU_1966 in out fe_tanh Vc=0.24886608795959314 Qo=8.774796100471918e-14 K=2.62 tau=9.967989058571382e-08 off=-0.2

*Grain_1967:
XU_1967 in out fe_tanh Vc=0.16706687154232475 Qo=5.89062875117664e-14 K=2.62 tau=1.0273718796081063e-07 off=-0.2

*Grain_1968:
XU_1968 in out fe_tanh Vc=0.2777013164342145 Qo=9.791500515484082e-14 K=2.62 tau=8.765752420080102e-08 off=-0.2

*Grain_1969:
XU_1969 in out fe_tanh Vc=0.2272364626083933 Qo=8.012154819201034e-14 K=2.62 tau=1.0559353648751127e-07 off=-0.2

*Grain_1970:
XU_1970 in out fe_tanh Vc=0.7944151214174554 Qo=2.801036801246148e-13 K=2.62 tau=9.795266510314351e-08 off=-0.2

*Grain_1971:
XU_1971 in out fe_tanh Vc=0.37724984832177527 Qo=1.3301492883574429e-13 K=2.62 tau=1.1306982452044215e-07 off=-0.2

*Grain_1972:
XU_1972 in out fe_tanh Vc=-0.1775050238914147 Qo=6.25866868494133e-14 K=2.62 tau=1.0210848922068196e-07 off=-0.2

*Grain_1973:
XU_1973 in out fe_tanh Vc=-0.011494391572845486 Qo=4.052819858970822e-15 K=2.62 tau=9.128109886843875e-08 off=-0.2

*Grain_1974:
XU_1974 in out fe_tanh Vc=0.5951353770630357 Qo=2.0983942122132387e-13 K=2.62 tau=1.1133643390761287e-07 off=-0.2

*Grain_1975:
XU_1975 in out fe_tanh Vc=-0.04018092901225834 Qo=1.4167436877432234e-14 K=2.62 tau=1.0787736103520611e-07 off=-0.2

*Grain_1976:
XU_1976 in out fe_tanh Vc=0.5076403269970505 Qo=1.7898944763013465e-13 K=2.62 tau=8.863866914351787e-08 off=-0.2

*Grain_1977:
XU_1977 in out fe_tanh Vc=0.5043649495424947 Qo=1.778345787787194e-13 K=2.62 tau=1.0561099265072679e-07 off=-0.2

*Grain_1978:
XU_1978 in out fe_tanh Vc=0.8987041175963711 Qo=3.168750491968631e-13 K=2.62 tau=1.0019550156734069e-07 off=-0.2

*Grain_1979:
XU_1979 in out fe_tanh Vc=0.5617777296486642 Qo=1.9807781252435795e-13 K=2.62 tau=9.158816305557853e-08 off=-0.2

*Grain_1980:
XU_1980 in out fe_tanh Vc=0.9291990039228166 Qo=3.2762727388989053e-13 K=2.62 tau=1.0164586542861982e-07 off=-0.2

*Grain_1981:
XU_1981 in out fe_tanh Vc=0.8222988186801544 Qo=2.8993522286366394e-13 K=2.62 tau=8.848630437123393e-08 off=-0.2

*Grain_1982:
XU_1982 in out fe_tanh Vc=0.5653593502951693 Qo=1.9934065999144331e-13 K=2.62 tau=8.988670502391775e-08 off=-0.2

*Grain_1983:
XU_1983 in out fe_tanh Vc=0.4440822513431344 Qo=1.5657943753297613e-13 K=2.62 tau=9.379232233402285e-08 off=-0.2

*Grain_1984:
XU_1984 in out fe_tanh Vc=0.79145192557564 Qo=2.7905888372302884e-13 K=2.62 tau=1.0572278355808962e-07 off=-0.2

*Grain_1985:
XU_1985 in out fe_tanh Vc=0.1532486185256568 Qo=5.4034094852649295e-14 K=2.62 tau=1.1375144365501483e-07 off=-0.2

*Grain_1986:
XU_1986 in out fe_tanh Vc=0.13731986466164225 Qo=4.841775843504844e-14 K=2.62 tau=8.862610036115062e-08 off=-0.2

*Grain_1987:
XU_1987 in out fe_tanh Vc=0.20760161482062453 Qo=7.31984761409301e-14 K=2.62 tau=1.0410826496754692e-07 off=-0.2

*Grain_1988:
XU_1988 in out fe_tanh Vc=-0.09836101974066752 Qo=3.4681217498745215e-14 K=2.62 tau=1.1021041062993914e-07 off=-0.2

*Grain_1989:
XU_1989 in out fe_tanh Vc=0.46228576513301106 Qo=1.629978339938162e-13 K=2.62 tau=1.0089509376234582e-07 off=-0.2

*Grain_1990:
XU_1990 in out fe_tanh Vc=0.13037855158629869 Qo=4.59703134092895e-14 K=2.62 tau=8.884286693080087e-08 off=-0.2

*Grain_1991:
XU_1991 in out fe_tanh Vc=0.2937404026668562 Qo=1.0357024378069042e-13 K=2.62 tau=9.273419001315554e-08 off=-0.2

*Grain_1992:
XU_1992 in out fe_tanh Vc=0.31919056047149497 Qo=1.1254374223086088e-13 K=2.62 tau=1.1176423518709599e-07 off=-0.2

*Grain_1993:
XU_1993 in out fe_tanh Vc=0.8180024399481405 Qo=2.8842035807622264e-13 K=2.62 tau=9.509451588828706e-08 off=-0.2

*Grain_1994:
XU_1994 in out fe_tanh Vc=0.31823067782216374 Qo=1.122052961775107e-13 K=2.62 tau=9.002044657966129e-08 off=-0.2

*Grain_1995:
XU_1995 in out fe_tanh Vc=0.6955093650702916 Qo=2.4523039336124387e-13 K=2.62 tau=1.1256443043790048e-07 off=-0.2

*Grain_1996:
XU_1996 in out fe_tanh Vc=0.366079519520935 Qo=1.2907637061729722e-13 K=2.62 tau=1.1029190992328387e-07 off=-0.2

*Grain_1997:
XU_1997 in out fe_tanh Vc=0.24507588780086795 Qo=8.64115702635994e-14 K=2.62 tau=8.854655881072479e-08 off=-0.2

*Grain_1998:
XU_1998 in out fe_tanh Vc=0.1432305570870831 Qo=5.050181581992879e-14 K=2.62 tau=1.0777103480374031e-07 off=-0.2

*Grain_1999:
XU_1999 in out fe_tanh Vc=0.43073812103283743 Qo=1.5187441630766583e-13 K=2.62 tau=1.0797173304491189e-07 off=-0.2
Rp in out R=50000.0
Cp in out 1.9e-10
.lib C:\Users\MBX\Desktop\Investigacion\Spice-LK-Model\Fe_model\fe_tanh.sp
.ends
